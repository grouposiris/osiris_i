// This is the unpowered netlist.
module core (clk,
    o_mem_write_M,
    rst,
    i_instr_ID,
    i_read_data_M,
    o_data_addr_M,
    o_funct3_MEM,
    o_pc_IF,
    o_write_data_M);
 input clk;
 output o_mem_write_M;
 input rst;
 input [31:0] i_instr_ID;
 input [31:0] i_read_data_M;
 output [31:0] o_data_addr_M;
 output [2:0] o_funct3_MEM;
 output [31:0] o_pc_IF;
 output [31:0] o_write_data_M;

 wire net469;
 wire net470;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ;
 wire \U_CONTROL_UNIT.i_branch_EX ;
 wire \U_CONTROL_UNIT.i_jump_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_mem_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_reg_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_reg_write_M ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.o_addr_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[9] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[10] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[11] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[12] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[13] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[14] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[15] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[16] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[17] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[18] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[19] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[20] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[21] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[22] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[23] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[24] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[25] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[26] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[27] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[28] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[29] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[2] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[30] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[31] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[3] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[4] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[5] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[6] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[7] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[8] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[9] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[11] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[19] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[24] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[25] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[26] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[27] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[28] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[29] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net47;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A (.DIODE(net2113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__B (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A_N (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__B (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__C (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A1 (.DIODE(net1655));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__C1 (.DIODE(\U_DATAPATH.U_EX_MEM.o_reg_write_M ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A0 (.DIODE(net2205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A2 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__B (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__C (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A1 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A1 (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A2 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A_N (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A_N (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__B (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__C (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__C (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A1 (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A2 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__B (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__C (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A1 (.DIODE(net1701));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A (.DIODE(net1701));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B2 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__C (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A_N (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__C (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__B1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1 (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A2 (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A_N (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__C (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A1 (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__B (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__C (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__B (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__C (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A2 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__B (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__C (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A1 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A2 (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__C (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A1 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A2 (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__B (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A_N (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__C (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(net2058));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A0 (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B1 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A0 (.DIODE(net2177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A1 (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__B1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__B (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__C (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A2 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A1 (.DIODE(net2023));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(net2023));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__B (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__S1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__C (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A2 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__C (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(net2125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A1 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A (.DIODE(net2125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(net2182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__C (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A0 (.DIODE(net2155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__B (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A2 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__C (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A_N (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A_N (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A1 (.DIODE(net2163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__B (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B2 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A1 (.DIODE(net2163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B2 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A3 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B1 (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A1 (.DIODE(net2103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A1 (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A2 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A1 (.DIODE(net2330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A2 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__C1 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A_N (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A1 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A_N (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A_N (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A2 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__B2 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A2 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A_N (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A_N (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A (.DIODE(net2155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(net2155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A (.DIODE(net2113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(net2113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A (.DIODE(net2177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A (.DIODE(net2177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__B (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A (.DIODE(net2205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A (.DIODE(net2205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__B (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__B (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A1 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A2 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__B (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A2 (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__S (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__S (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__S (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A1 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A1 (.DIODE(net2028));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__S (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A1 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A0 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(net2043));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A1 (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__S (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A0 (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(_1936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__S (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A0 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__S (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A (.DIODE(_1936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__C (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__B (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__B (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__S (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A2 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__B (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A2 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A1 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A2 (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A0 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(net2043));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B1 (.DIODE(_1936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__D (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__B (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__D_N (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__D (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__C_N (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__B (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A (.DIODE(net2106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__B (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A (.DIODE(net2056));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(net2221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__B (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A (.DIODE(net2095));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__B (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__C (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A1 (.DIODE(net1959));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__C (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(net2106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__C (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A (.DIODE(net2056));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A1 (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B2 (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(net2042));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B2 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A1 (.DIODE(net1959));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__B2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__B (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__D_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__D_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__B (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__B (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__D_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B2 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A3 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A1 (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__C (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A3 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__C (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__C (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__C (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A3 (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__D (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__C (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A3 (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A3 (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__C1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A (.DIODE(net1701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A (.DIODE(net1655));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A (.DIODE(net2023));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A (.DIODE(net2058));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A (.DIODE(net2103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__B (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(net2125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A (.DIODE(net2163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__B (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B (.DIODE(net2182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A0 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A0 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__C1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A0 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A0 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A1 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A0 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A0 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A0 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A1 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A0 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A0 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A0 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A1 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__C (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__C (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__C1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A0 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__S1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A0 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A0 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A0 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A3 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__C (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B2 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A3 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__S0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A0 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A3 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__S0 (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__S1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A0 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A3 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__S0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A0 (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__S (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__B1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1_N (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B1 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A2 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A0 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A0 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A3 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A3 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__S (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A2 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A2 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A3 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A0 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A3 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__S1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A2 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B1 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__C1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A0 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A1 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A2 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__S1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__B2 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__C1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A0 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__S (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A0 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__B1_N (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A2 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A0 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A1 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A3 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__S0 (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__S1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__B1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__B2 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A2 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A2 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A1 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A0 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A3 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B2 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A2 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A0 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A1 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1_N (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__B2 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A1 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__B1 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A2 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A0 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A2 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A3 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__S1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__B1_N (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A2 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__C1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A1 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__B1_N (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__S (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A2 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A0 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A2 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A3 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A1 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A2 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__C1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__B1_N (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A0 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__S (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A2 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__B1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A0 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A2 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A3 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__S1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__B1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A2 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A1 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A0 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A2 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A3 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__S0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__B1_N (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A2 (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A0 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A1_N (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A2_N (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__B1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__B2 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__B (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__C1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A3 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A1_N (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A2 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A3 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B1 (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A1 (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A1 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A0 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A1 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A2 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__C1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A1_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A0 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A2 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A3 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__S1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B1 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B2 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A0 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B1 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__B2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A0 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A3 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A1_N (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__B1 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__C1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A0 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1_N (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__B1 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__B1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A2 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A0 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A3 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__S1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A1_N (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__B1 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A1 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A1 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__B1 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A3 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A1 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__B1 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__B2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__B1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__C1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A2 (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__B1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__B (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A (.DIODE(net1959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A (.DIODE(net2042));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A (.DIODE(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A (.DIODE(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A (.DIODE(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(net2126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__C1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__C (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A2 (.DIODE(_3447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A2 (.DIODE(_3447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A1 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A1 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A1 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A1 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A (.DIODE(net1959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A (.DIODE(net2042));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A (.DIODE(net2221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A (.DIODE(net2056));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A (.DIODE(net2106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__S (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A1 (.DIODE(net2043));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A1 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__D (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__SET_B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__D (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__D (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7562__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__D (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__D (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__CLK (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__D (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7566__D (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__D (.DIODE(_0594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__D (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__D (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__D (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__D (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__D (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__D (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__D (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8286__D (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(_3457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(_3457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(_3455_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(_3455_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(_3453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(_3453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(_3447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(_3435_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(_3435_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(_3451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(_3451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(net2054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(net2054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout396_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout399_A (.DIODE(net2126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(net2233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net2233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(net2233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(net2263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(net2263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(net2095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout444_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout445_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout449_A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout450_A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1160_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1168_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1175_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1222_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1275_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1412_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1430_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1437_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1467_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1468_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1469_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1477_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1478_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1482_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1518_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1528_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1529_A (.DIODE(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1535_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1536_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1539_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1540_A (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1549_A (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1550_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1556_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1567_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1590_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1597_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1606_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1607_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1610_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1611_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1614_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1627_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1629_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1633_A (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1650_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1651_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1656_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1658_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1662_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1669_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1673_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1674_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1680_A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1684_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1685_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1687_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1696_A (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1698_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1704_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1709_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1721_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1727_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1730_A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1746_A (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1753_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1760_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1766_A (.DIODE(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1767_A (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1771_A (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1772_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1777_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1785_A (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1787_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1791_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1794_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1795_A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1798_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1806_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1807_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1810_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1812_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1814_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1816_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1819_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1822_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1823_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1824_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1827_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1830_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1833_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1836_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1837_A (.DIODE(\U_DATAPATH.U_EX_MEM.o_reg_write_M ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1840_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1842_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1843_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1844_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1847_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1848_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1850_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1851_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1852_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold384_A (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold498_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3572_ (.A(net578),
    .Y(_1277_));
 sky130_fd_sc_hd__inv_2 _3573_ (.A(net2119),
    .Y(_1278_));
 sky130_fd_sc_hd__inv_2 _3574_ (.A(net2148),
    .Y(_1279_));
 sky130_fd_sc_hd__inv_2 _3575_ (.A(net2170),
    .Y(_1280_));
 sky130_fd_sc_hd__inv_2 _3576_ (.A(net2029),
    .Y(_1281_));
 sky130_fd_sc_hd__inv_2 _3577_ (.A(net2037),
    .Y(_1282_));
 sky130_fd_sc_hd__inv_2 _3578_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1283_));
 sky130_fd_sc_hd__inv_2 _3579_ (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .Y(_1284_));
 sky130_fd_sc_hd__inv_2 _3580_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .Y(_1285_));
 sky130_fd_sc_hd__inv_2 _3581_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_1286_));
 sky130_fd_sc_hd__inv_2 _3582_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1287_));
 sky130_fd_sc_hd__inv_2 _3583_ (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .Y(_1288_));
 sky130_fd_sc_hd__inv_2 _3584_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .Y(_1289_));
 sky130_fd_sc_hd__inv_2 _3585_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .Y(_1290_));
 sky130_fd_sc_hd__inv_2 _3586_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .Y(_1291_));
 sky130_fd_sc_hd__inv_2 _3587_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .Y(_1292_));
 sky130_fd_sc_hd__inv_2 _3588_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .Y(_1293_));
 sky130_fd_sc_hd__inv_2 _3589_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .Y(_1294_));
 sky130_fd_sc_hd__inv_2 _3590_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _3591_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .Y(_1296_));
 sky130_fd_sc_hd__inv_2 _3592_ (.A(net2113),
    .Y(_1297_));
 sky130_fd_sc_hd__inv_2 _3593_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .Y(_1298_));
 sky130_fd_sc_hd__inv_2 _3594_ (.A(net2306),
    .Y(_1299_));
 sky130_fd_sc_hd__inv_2 _3595_ (.A(net2290),
    .Y(_1300_));
 sky130_fd_sc_hd__inv_2 _3596_ (.A(net2045),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_6 _3597_ (.A(net457),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _3598__1 (.A(clknet_leaf_36_clk),
    .Y(net473));
 sky130_fd_sc_hd__or2_1 _3599_ (.A(net385),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_1302_));
 sky130_fd_sc_hd__nand2_1 _3600_ (.A(net385),
    .B(net2059),
    .Y(_1303_));
 sky130_fd_sc_hd__or2_1 _3601_ (.A(net395),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_1304_));
 sky130_fd_sc_hd__nand2_1 _3602_ (.A(net395),
    .B(net2006),
    .Y(_1305_));
 sky130_fd_sc_hd__a22o_1 _3603_ (.A1(_1302_),
    .A2(_1303_),
    .B1(_1304_),
    .B2(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__or2_1 _3604_ (.A(net369),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_1 _3605_ (.A(net369),
    .B(net1631),
    .Y(_1308_));
 sky130_fd_sc_hd__or2_1 _3606_ (.A(net374),
    .B(net2167),
    .X(_1309_));
 sky130_fd_sc_hd__nand2_1 _3607_ (.A(net374),
    .B(net1308),
    .Y(_1310_));
 sky130_fd_sc_hd__a22o_1 _3608_ (.A1(_1307_),
    .A2(_1308_),
    .B1(_1309_),
    .B2(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__or2_1 _3609_ (.A(net423),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_1312_));
 sky130_fd_sc_hd__nand2_1 _3610_ (.A(net423),
    .B(net2006),
    .Y(_1313_));
 sky130_fd_sc_hd__or2_1 _3611_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_1314_));
 sky130_fd_sc_hd__nand2_1 _3612_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .B(net1631),
    .Y(_1315_));
 sky130_fd_sc_hd__or2_1 _3613_ (.A(net414),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_1316_));
 sky130_fd_sc_hd__nand2_1 _3614_ (.A(net414),
    .B(net2059),
    .Y(_1317_));
 sky130_fd_sc_hd__or2_1 _3615_ (.A(net403),
    .B(net2167),
    .X(_1318_));
 sky130_fd_sc_hd__nand2_1 _3616_ (.A(net403),
    .B(net1308),
    .Y(_1319_));
 sky130_fd_sc_hd__a22o_1 _3617_ (.A1(_1312_),
    .A2(_1313_),
    .B1(_1316_),
    .B2(_1317_),
    .X(_1320_));
 sky130_fd_sc_hd__a22o_1 _3618_ (.A1(_1314_),
    .A2(_1315_),
    .B1(_1318_),
    .B2(_1319_),
    .X(_1321_));
 sky130_fd_sc_hd__o22a_2 _3619_ (.A1(_1306_),
    .A2(_1311_),
    .B1(_1320_),
    .B2(net2168),
    .X(_1322_));
 sky130_fd_sc_hd__nor3b_4 _3620_ (.A(net1282),
    .B(_1322_),
    .C_N(net1619),
    .Y(_1323_));
 sky130_fd_sc_hd__or3b_4 _3621_ (.A(net1282),
    .B(net2169),
    .C_N(net1619),
    .X(_1324_));
 sky130_fd_sc_hd__nand2b_1 _3622_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1325_));
 sky130_fd_sc_hd__and2b_1 _3623_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1326_));
 sky130_fd_sc_hd__nand2b_1 _3624_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1327_));
 sky130_fd_sc_hd__nor4_1 _3625_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1328_));
 sky130_fd_sc_hd__a221o_1 _3626_ (.A1(_1283_),
    .A2(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B1(_1284_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .C1(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__nand2_1 _3627_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1330_));
 sky130_fd_sc_hd__or2_1 _3628_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(_1331_));
 sky130_fd_sc_hd__a21o_1 _3629_ (.A1(_1330_),
    .A2(_1331_),
    .B1(_1328_),
    .X(_1332_));
 sky130_fd_sc_hd__o2111ai_4 _3630_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .A2(_1284_),
    .B1(_1325_),
    .C1(_1327_),
    .D1(net851),
    .Y(_1333_));
 sky130_fd_sc_hd__nor3_4 _3631_ (.A(_1329_),
    .B(_1332_),
    .C(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__or3_4 _3632_ (.A(_1329_),
    .B(_1332_),
    .C(_1333_),
    .X(_1335_));
 sky130_fd_sc_hd__nand2b_1 _3633_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2b_1 _3634_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2b_1 _3635_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_1339_));
 sky130_fd_sc_hd__or2_1 _3637_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_1340_));
 sky130_fd_sc_hd__a21oi_1 _3638_ (.A1(_1339_),
    .A2(_1340_),
    .B1(_1328_),
    .Y(_1341_));
 sky130_fd_sc_hd__o221a_1 _3639_ (.A1(_1283_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B1(_1286_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .C1(_1337_),
    .X(_1342_));
 sky130_fd_sc_hd__o2111a_1 _3640_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .A2(_1285_),
    .B1(_1336_),
    .C1(_1338_),
    .D1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1343_));
 sky130_fd_sc_hd__and3_4 _3641_ (.A(_1341_),
    .B(_1342_),
    .C(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__and2_4 _3642_ (.A(net303),
    .B(net302),
    .X(_1345_));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(net364),
    .B(net366),
    .Y(_1346_));
 sky130_fd_sc_hd__and2b_1 _3644_ (.A_N(net366),
    .B(net364),
    .X(_1347_));
 sky130_fd_sc_hd__and2_1 _3645_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .X(_1348_));
 sky130_fd_sc_hd__mux4_2 _3646_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ),
    .A1(net34),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ),
    .S0(net364),
    .S1(net366),
    .X(_1349_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__and3_1 _3648_ (.A(net303),
    .B(net302),
    .C(_1349_),
    .X(_1351_));
 sky130_fd_sc_hd__nor2_2 _3649_ (.A(net304),
    .B(_1344_),
    .Y(_1352_));
 sky130_fd_sc_hd__a221o_2 _3650_ (.A1(net1655),
    .A2(_1334_),
    .B1(net242),
    .B2(net2269),
    .C1(_1351_),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_4 _3651_ (.A0(net2098),
    .A1(_1353_),
    .S(net362),
    .X(_1354_));
 sky130_fd_sc_hd__or4_1 _3652_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .X(_1355_));
 sky130_fd_sc_hd__o2bb2a_4 _3653_ (.A1_N(_1292_),
    .A2_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B1(_1284_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1356_));
 sky130_fd_sc_hd__o22a_1 _3654_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .A2(_1291_),
    .B1(_1292_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1357_));
 sky130_fd_sc_hd__a22oi_2 _3655_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1290_),
    .B1(_1291_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1358_));
 sky130_fd_sc_hd__o211a_1 _3656_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1290_),
    .B1(_1355_),
    .C1(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(_1359_));
 sky130_fd_sc_hd__o2111a_4 _3657_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .A2(_1289_),
    .B1(_1357_),
    .C1(_1358_),
    .D1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__and2_1 _3658_ (.A(net332),
    .B(net301),
    .X(_1361_));
 sky130_fd_sc_hd__and2b_1 _3659_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1362_));
 sky130_fd_sc_hd__a221o_1 _3660_ (.A1(_1285_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .B1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .B2(_1287_),
    .C1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__xor2_1 _3661_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _3662_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .A2(_1290_),
    .B1(_1292_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__o211a_1 _3663_ (.A1(_1286_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B1(_1355_),
    .C1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1366_));
 sky130_fd_sc_hd__or3b_2 _3664_ (.A(_1363_),
    .B(_1365_),
    .C_N(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__a21oi_4 _3665_ (.A1(net331),
    .A2(net300),
    .B1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__and3_1 _3666_ (.A(net67),
    .B(net331),
    .C(net300),
    .X(_1369_));
 sky130_fd_sc_hd__a21boi_4 _3667_ (.A1(net331),
    .A2(net300),
    .B1_N(_1367_),
    .Y(_1370_));
 sky130_fd_sc_hd__a221o_4 _3668_ (.A1(_1349_),
    .A2(net241),
    .B1(net239),
    .B2(net2329),
    .C1(_1369_),
    .X(_1371_));
 sky130_fd_sc_hd__inv_2 _3669_ (.A(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__xnor2_1 _3670_ (.A(_1354_),
    .B(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__mux4_2 _3671_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ),
    .A1(net33),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ),
    .S0(net365),
    .S1(net367),
    .X(_1374_));
 sky130_fd_sc_hd__a22o_1 _3672_ (.A1(net2201),
    .A2(net242),
    .B1(_1374_),
    .B2(_1345_),
    .X(_1375_));
 sky130_fd_sc_hd__a21oi_4 _3673_ (.A1(net2166),
    .A2(net305),
    .B1(net2202),
    .Y(_1376_));
 sky130_fd_sc_hd__inv_2 _3674_ (.A(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux2_2 _3675_ (.A0(_1295_),
    .A1(_1376_),
    .S(net362),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _3676_ (.A0(net2205),
    .A1(_1377_),
    .S(net362),
    .X(_1379_));
 sky130_fd_sc_hd__and3_1 _3677_ (.A(net66),
    .B(net332),
    .C(net301),
    .X(_1380_));
 sky130_fd_sc_hd__a221o_4 _3678_ (.A1(net2308),
    .A2(net238),
    .B1(net361),
    .B2(net240),
    .C1(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__a21oi_1 _3679_ (.A1(_1378_),
    .A2(_1381_),
    .B1(_1373_),
    .Y(_1382_));
 sky130_fd_sc_hd__nor2_1 _3680_ (.A(_1378_),
    .B(_1381_),
    .Y(_1383_));
 sky130_fd_sc_hd__mux4_2 _3681_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ),
    .A1(net35),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ),
    .S0(net365),
    .S1(net367),
    .X(_1384_));
 sky130_fd_sc_hd__and3_1 _3682_ (.A(net303),
    .B(net302),
    .C(net360),
    .X(_1385_));
 sky130_fd_sc_hd__a221o_2 _3683_ (.A1(net2187),
    .A2(net305),
    .B1(net242),
    .B2(net2268),
    .C1(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_2 _3684_ (.A0(net2171),
    .A1(_1386_),
    .S(net363),
    .X(_1387_));
 sky130_fd_sc_hd__and3_1 _3685_ (.A(net68),
    .B(net332),
    .C(net301),
    .X(_1388_));
 sky130_fd_sc_hd__a221o_4 _3686_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .A2(net238),
    .B1(net360),
    .B2(net240),
    .C1(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__inv_2 _3687_ (.A(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__and2_1 _3688_ (.A(_1387_),
    .B(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__mux4_2 _3689_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ),
    .A1(net62),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ),
    .S0(net364),
    .S1(net366),
    .X(_1392_));
 sky130_fd_sc_hd__a22o_1 _3690_ (.A1(net2084),
    .A2(net243),
    .B1(net359),
    .B2(_1345_),
    .X(_1393_));
 sky130_fd_sc_hd__a21oi_4 _3691_ (.A1(net860),
    .A2(_1334_),
    .B1(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2_1 _3692_ (.A(net2302),
    .B(net2215),
    .Y(_1395_));
 sky130_fd_sc_hd__o21ai_4 _3693_ (.A1(net2302),
    .A2(_1394_),
    .B1(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__and3_1 _3694_ (.A(net95),
    .B(net331),
    .C(net300),
    .X(_1397_));
 sky130_fd_sc_hd__a221o_4 _3695_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .A2(net239),
    .B1(net359),
    .B2(net241),
    .C1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__and2b_1 _3696_ (.A_N(_1398_),
    .B(_1396_),
    .X(_1399_));
 sky130_fd_sc_hd__nand2b_1 _3697_ (.A_N(_1396_),
    .B(_1398_),
    .Y(_1400_));
 sky130_fd_sc_hd__or4b_1 _3698_ (.A(_1383_),
    .B(_1391_),
    .C(_1399_),
    .D_N(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__mux4_2 _3699_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ),
    .A1(net61),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ),
    .S0(net364),
    .S1(net366),
    .X(_1402_));
 sky130_fd_sc_hd__and3_1 _3700_ (.A(net303),
    .B(net302),
    .C(net358),
    .X(_1403_));
 sky130_fd_sc_hd__a221o_2 _3701_ (.A1(net2192),
    .A2(net305),
    .B1(net242),
    .B2(net2281),
    .C1(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_2 _3702_ (.A0(net2138),
    .A1(_1404_),
    .S(net363),
    .X(_1405_));
 sky130_fd_sc_hd__and3_1 _3703_ (.A(net2192),
    .B(net331),
    .C(net300),
    .X(_1406_));
 sky130_fd_sc_hd__a221o_4 _3704_ (.A1(net2315),
    .A2(net239),
    .B1(net358),
    .B2(net241),
    .C1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__and2b_1 _3705_ (.A_N(_1407_),
    .B(_1405_),
    .X(_1408_));
 sky130_fd_sc_hd__and2b_1 _3706_ (.A_N(_1405_),
    .B(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__or2_1 _3707_ (.A(_1408_),
    .B(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__inv_2 _3708_ (.A(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux4_2 _3709_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ),
    .A1(net32),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ),
    .S0(net365),
    .S1(net367),
    .X(_1412_));
 sky130_fd_sc_hd__and3_1 _3710_ (.A(net303),
    .B(net302),
    .C(net357),
    .X(_1413_));
 sky130_fd_sc_hd__a221o_2 _3711_ (.A1(net2087),
    .A2(net305),
    .B1(net242),
    .B2(net2132),
    .C1(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_2 _3712_ (.A0(net2211),
    .A1(_1414_),
    .S(net363),
    .X(_1415_));
 sky130_fd_sc_hd__and3_1 _3713_ (.A(net2087),
    .B(net332),
    .C(net301),
    .X(_1416_));
 sky130_fd_sc_hd__a221o_4 _3714_ (.A1(net2316),
    .A2(net238),
    .B1(net357),
    .B2(net240),
    .C1(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__xnor2_1 _3715_ (.A(_1415_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__and4b_1 _3716_ (.A_N(_1401_),
    .B(_1418_),
    .C(_1411_),
    .D(_1382_),
    .X(_1419_));
 sky130_fd_sc_hd__mux4_2 _3717_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ),
    .A1(net57),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ),
    .S0(net364),
    .S1(net366),
    .X(_1420_));
 sky130_fd_sc_hd__and2_1 _3718_ (.A(net1007),
    .B(net304),
    .X(_1421_));
 sky130_fd_sc_hd__a221oi_4 _3719_ (.A1(net2222),
    .A2(net243),
    .B1(net356),
    .B2(_1345_),
    .C1(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__nand2_1 _3720_ (.A(net2302),
    .B(net2273),
    .Y(_1423_));
 sky130_fd_sc_hd__mux2_1 _3721_ (.A0(_1294_),
    .A1(_1422_),
    .S(net363),
    .X(_1424_));
 sky130_fd_sc_hd__o21ai_4 _3722_ (.A1(net2302),
    .A2(_1422_),
    .B1(_1423_),
    .Y(_1425_));
 sky130_fd_sc_hd__and3_1 _3723_ (.A(net1007),
    .B(net331),
    .C(net300),
    .X(_1426_));
 sky130_fd_sc_hd__a221o_4 _3724_ (.A1(net2343),
    .A2(net239),
    .B1(net356),
    .B2(net241),
    .C1(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(net214),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__or2_1 _3726_ (.A(net214),
    .B(_1427_),
    .X(_1429_));
 sky130_fd_sc_hd__mux4_2 _3727_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ),
    .A1(net56),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ),
    .S0(net364),
    .S1(net366),
    .X(_1430_));
 sky130_fd_sc_hd__and3_1 _3728_ (.A(net303),
    .B(net302),
    .C(net355),
    .X(_1431_));
 sky130_fd_sc_hd__a221oi_4 _3729_ (.A1(net1701),
    .A2(net304),
    .B1(net243),
    .B2(net2193),
    .C1(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__inv_2 _3730_ (.A(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__mux2_1 _3731_ (.A0(_1293_),
    .A1(_1432_),
    .S(net363),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_2 _3732_ (.A0(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .A1(_1433_),
    .S(net363),
    .X(_1435_));
 sky130_fd_sc_hd__and3_1 _3733_ (.A(net1701),
    .B(net331),
    .C(net300),
    .X(_1436_));
 sky130_fd_sc_hd__a221o_4 _3734_ (.A1(net2328),
    .A2(net239),
    .B1(net355),
    .B2(net241),
    .C1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__a22oi_2 _3735_ (.A1(_1428_),
    .A2(_1429_),
    .B1(net210),
    .B2(_1437_),
    .Y(_1438_));
 sky130_fd_sc_hd__a22o_1 _3736_ (.A1(net42),
    .A2(_1347_),
    .B1(_1348_),
    .B2(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ),
    .X(_1439_));
 sky130_fd_sc_hd__a21o_1 _3737_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ),
    .A2(_1346_),
    .B1(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__and3_1 _3738_ (.A(net2086),
    .B(net331),
    .C(net300),
    .X(_1441_));
 sky130_fd_sc_hd__a221o_2 _3739_ (.A1(net2301),
    .A2(net239),
    .B1(net299),
    .B2(net241),
    .C1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__inv_2 _3740_ (.A(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__and3_1 _3741_ (.A(net303),
    .B(net302),
    .C(net299),
    .X(_1444_));
 sky130_fd_sc_hd__and2_1 _3742_ (.A(net2086),
    .B(net304),
    .X(_1445_));
 sky130_fd_sc_hd__and3b_2 _3743_ (.A_N(_1344_),
    .B(net2336),
    .C(_1335_),
    .X(_1446_));
 sky130_fd_sc_hd__o31ai_2 _3744_ (.A1(_1444_),
    .A2(_1445_),
    .A3(_1446_),
    .B1(net363),
    .Y(_1447_));
 sky130_fd_sc_hd__nand2_1 _3745_ (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .B(net826),
    .Y(_1448_));
 sky130_fd_sc_hd__and2_2 _3746_ (.A(_1447_),
    .B(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_1 _3747_ (.A(_1447_),
    .B(_1448_),
    .Y(_1450_));
 sky130_fd_sc_hd__xnor2_1 _3748_ (.A(_1443_),
    .B(net206),
    .Y(_1451_));
 sky130_fd_sc_hd__nor2_1 _3749_ (.A(net210),
    .B(_1437_),
    .Y(_1452_));
 sky130_fd_sc_hd__mux4_2 _3750_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ),
    .A1(net58),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ),
    .S0(net364),
    .S1(net366),
    .X(_1453_));
 sky130_fd_sc_hd__a22o_1 _3751_ (.A1(net2164),
    .A2(net243),
    .B1(net354),
    .B2(_1345_),
    .X(_1454_));
 sky130_fd_sc_hd__a21oi_4 _3752_ (.A1(net2100),
    .A2(net304),
    .B1(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _3753_ (.A(net2302),
    .B(net2067),
    .Y(_1456_));
 sky130_fd_sc_hd__o21ai_4 _3754_ (.A1(net2302),
    .A2(_1455_),
    .B1(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__and3_1 _3755_ (.A(net91),
    .B(net331),
    .C(net300),
    .X(_1458_));
 sky130_fd_sc_hd__a221o_4 _3756_ (.A1(net2311),
    .A2(net239),
    .B1(net354),
    .B2(net241),
    .C1(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__and2b_1 _3757_ (.A_N(_1459_),
    .B(_1457_),
    .X(_1460_));
 sky130_fd_sc_hd__nor2_1 _3758_ (.A(_1452_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__mux4_1 _3759_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ),
    .A1(net53),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ),
    .S0(net364),
    .S1(net366),
    .X(_1462_));
 sky130_fd_sc_hd__and3_1 _3760_ (.A(_1335_),
    .B(_1344_),
    .C(net353),
    .X(_1463_));
 sky130_fd_sc_hd__a221oi_4 _3761_ (.A1(net86),
    .A2(net304),
    .B1(net243),
    .B2(net2344),
    .C1(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .B(net2226),
    .Y(_1465_));
 sky130_fd_sc_hd__o21a_1 _3763_ (.A1(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .A2(_1464_),
    .B1(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__o21ai_4 _3764_ (.A1(net2302),
    .A2(_1464_),
    .B1(_1465_),
    .Y(_1467_));
 sky130_fd_sc_hd__and3_1 _3765_ (.A(net86),
    .B(_1356_),
    .C(_1360_),
    .X(_1468_));
 sky130_fd_sc_hd__a221o_4 _3766_ (.A1(net2337),
    .A2(net239),
    .B1(net353),
    .B2(net241),
    .C1(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__xnor2_1 _3767_ (.A(_1467_),
    .B(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__a22o_1 _3768_ (.A1(net31),
    .A2(_1347_),
    .B1(_1348_),
    .B2(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ),
    .X(_1471_));
 sky130_fd_sc_hd__a21o_1 _3769_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ),
    .A2(_1346_),
    .B1(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__and3_1 _3770_ (.A(net303),
    .B(net302),
    .C(net298),
    .X(_1473_));
 sky130_fd_sc_hd__a221oi_4 _3771_ (.A1(net2129),
    .A2(net304),
    .B1(net243),
    .B2(net2291),
    .C1(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(net773),
    .B(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .Y(_1475_));
 sky130_fd_sc_hd__o21ai_4 _3773_ (.A1(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .A2(_1474_),
    .B1(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__and3_1 _3774_ (.A(net2129),
    .B(net331),
    .C(net300),
    .X(_1477_));
 sky130_fd_sc_hd__a221o_2 _3775_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .A2(net239),
    .B1(net298),
    .B2(net241),
    .C1(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__nand2_1 _3776_ (.A(net194),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__or2_1 _3777_ (.A(net194),
    .B(_1478_),
    .X(_1480_));
 sky130_fd_sc_hd__nand2_1 _3778_ (.A(_1479_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__and4_1 _3779_ (.A(_1451_),
    .B(_1461_),
    .C(_1470_),
    .D(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__mux4_2 _3780_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ),
    .A1(net59),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ),
    .S0(net364),
    .S1(net366),
    .X(_1483_));
 sky130_fd_sc_hd__and3_1 _3781_ (.A(_1335_),
    .B(_1344_),
    .C(net352),
    .X(_1484_));
 sky130_fd_sc_hd__a221o_2 _3782_ (.A1(net2146),
    .A2(net304),
    .B1(net243),
    .B2(net2261),
    .C1(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_2 _3783_ (.A0(net2235),
    .A1(_1485_),
    .S(net363),
    .X(_1486_));
 sky130_fd_sc_hd__and3_1 _3784_ (.A(net92),
    .B(net331),
    .C(net300),
    .X(_1487_));
 sky130_fd_sc_hd__a221o_4 _3785_ (.A1(net2265),
    .A2(_1370_),
    .B1(_1483_),
    .B2(net241),
    .C1(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__xor2_1 _3786_ (.A(_1486_),
    .B(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__mux4_2 _3787_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ),
    .A1(net60),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ),
    .S0(net364),
    .S1(net366),
    .X(_1490_));
 sky130_fd_sc_hd__and3_1 _3788_ (.A(net303),
    .B(net302),
    .C(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a221o_2 _3789_ (.A1(net2210),
    .A2(net304),
    .B1(net243),
    .B2(net2231),
    .C1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_2 _3790_ (.A0(net2188),
    .A1(_1492_),
    .S(net363),
    .X(_1493_));
 sky130_fd_sc_hd__and3_1 _3791_ (.A(net2210),
    .B(net331),
    .C(net300),
    .X(_1494_));
 sky130_fd_sc_hd__a221o_4 _3792_ (.A1(net2309),
    .A2(net239),
    .B1(net351),
    .B2(net241),
    .C1(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__or2_1 _3794_ (.A(_1493_),
    .B(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__nand2b_1 _3795_ (.A_N(_1457_),
    .B(_1459_),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_1 _3796_ (.A(_1493_),
    .B(_1496_),
    .Y(_1499_));
 sky130_fd_sc_hd__and4b_1 _3797_ (.A_N(_1489_),
    .B(_1497_),
    .C(_1498_),
    .D(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__mux4_2 _3798_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ),
    .A1(net36),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ),
    .S0(net364),
    .S1(net366),
    .X(_1501_));
 sky130_fd_sc_hd__and3_1 _3799_ (.A(_1335_),
    .B(_1344_),
    .C(net350),
    .X(_1502_));
 sky130_fd_sc_hd__a221o_4 _3800_ (.A1(net2133),
    .A2(net304),
    .B1(net243),
    .B2(net2278),
    .C1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_2 _3801_ (.A0(net2224),
    .A1(_1503_),
    .S(net363),
    .X(_1504_));
 sky130_fd_sc_hd__and3_1 _3802_ (.A(net69),
    .B(net331),
    .C(net300),
    .X(_1505_));
 sky130_fd_sc_hd__a221o_4 _3803_ (.A1(net2335),
    .A2(net239),
    .B1(net350),
    .B2(net241),
    .C1(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__xnor2_1 _3804_ (.A(_1504_),
    .B(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__mux4_2 _3805_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ),
    .A1(net37),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ),
    .S0(net364),
    .S1(net366),
    .X(_1508_));
 sky130_fd_sc_hd__and3_1 _3806_ (.A(_1335_),
    .B(_1344_),
    .C(net349),
    .X(_1509_));
 sky130_fd_sc_hd__a221o_1 _3807_ (.A1(net2092),
    .A2(net304),
    .B1(net243),
    .B2(net2197),
    .C1(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_2 _3808_ (.A0(net2088),
    .A1(_1510_),
    .S(net363),
    .X(_1511_));
 sky130_fd_sc_hd__and3_1 _3809_ (.A(net70),
    .B(net331),
    .C(net300),
    .X(_1512_));
 sky130_fd_sc_hd__a221o_4 _3810_ (.A1(net2325),
    .A2(_1370_),
    .B1(net349),
    .B2(net241),
    .C1(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2b_1 _3811_ (.A_N(_1511_),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__and2b_1 _3812_ (.A_N(_1513_),
    .B(_1511_),
    .X(_1515_));
 sky130_fd_sc_hd__inv_2 _3813_ (.A(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__o2111a_1 _3814_ (.A1(_1387_),
    .A2(_1390_),
    .B1(_1507_),
    .C1(_1514_),
    .D1(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__and4_1 _3815_ (.A(_1438_),
    .B(_1482_),
    .C(_1500_),
    .D(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__mux4_2 _3816_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ),
    .A1(net45),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ),
    .S0(net365),
    .S1(net367),
    .X(_1519_));
 sky130_fd_sc_hd__and3_1 _3817_ (.A(net303),
    .B(net302),
    .C(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__a221o_4 _3818_ (.A1(net2058),
    .A2(net304),
    .B1(net243),
    .B2(net2305),
    .C1(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_2 _3819_ (.A0(net2151),
    .A1(_1521_),
    .S(net362),
    .X(_1522_));
 sky130_fd_sc_hd__and3_1 _3820_ (.A(net78),
    .B(net332),
    .C(net301),
    .X(_1523_));
 sky130_fd_sc_hd__a221o_4 _3821_ (.A1(net2323),
    .A2(net238),
    .B1(net348),
    .B2(net240),
    .C1(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__xor2_1 _3822_ (.A(_1522_),
    .B(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__mux4_2 _3823_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ),
    .A1(net46),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ),
    .S0(net365),
    .S1(net367),
    .X(_1526_));
 sky130_fd_sc_hd__a22o_1 _3824_ (.A1(net2010),
    .A2(net242),
    .B1(_1526_),
    .B2(_1345_),
    .X(_1527_));
 sky130_fd_sc_hd__a21oi_4 _3825_ (.A1(net969),
    .A2(net305),
    .B1(net2011),
    .Y(_1528_));
 sky130_fd_sc_hd__inv_2 _3826_ (.A(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__mux2_2 _3827_ (.A0(_1298_),
    .A1(_1528_),
    .S(net362),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _3828_ (.A0(net2177),
    .A1(_1529_),
    .S(net362),
    .X(_1531_));
 sky130_fd_sc_hd__and3_1 _3829_ (.A(net969),
    .B(net332),
    .C(net301),
    .X(_1532_));
 sky130_fd_sc_hd__a221o_4 _3830_ (.A1(net2322),
    .A2(net238),
    .B1(net347),
    .B2(net240),
    .C1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__nor2_1 _3831_ (.A(_1530_),
    .B(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__mux4_2 _3832_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ),
    .A1(net44),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ),
    .S0(net365),
    .S1(net367),
    .X(_1535_));
 sky130_fd_sc_hd__a22o_1 _3833_ (.A1(net2249),
    .A2(net242),
    .B1(net346),
    .B2(_1345_),
    .X(_1536_));
 sky130_fd_sc_hd__a21oi_4 _3834_ (.A1(net2032),
    .A2(net305),
    .B1(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__inv_2 _3835_ (.A(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__mux2_2 _3836_ (.A0(net2077),
    .A1(_1538_),
    .S(net362),
    .X(_1539_));
 sky130_fd_sc_hd__and3_1 _3837_ (.A(net2032),
    .B(net332),
    .C(net301),
    .X(_1540_));
 sky130_fd_sc_hd__a221o_4 _3838_ (.A1(net2313),
    .A2(net238),
    .B1(net346),
    .B2(net240),
    .C1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__inv_2 _3839_ (.A(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__a2bb2o_1 _3840_ (.A1_N(_1542_),
    .A2_N(_1539_),
    .B1(_1533_),
    .B2(_1530_),
    .X(_1543_));
 sky130_fd_sc_hd__or3_2 _3841_ (.A(_1525_),
    .B(_1534_),
    .C(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__mux4_2 _3842_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ),
    .A1(net38),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ),
    .S0(net364),
    .S1(net366),
    .X(_1545_));
 sky130_fd_sc_hd__a22o_1 _3843_ (.A1(net2345),
    .A2(net243),
    .B1(net345),
    .B2(_1345_),
    .X(_1546_));
 sky130_fd_sc_hd__a21oi_4 _3844_ (.A1(net2223),
    .A2(net304),
    .B1(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__inv_2 _3845_ (.A(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__mux2_2 _3846_ (.A0(net2134),
    .A1(_1548_),
    .S(net363),
    .X(_1549_));
 sky130_fd_sc_hd__and3_1 _3847_ (.A(net71),
    .B(net331),
    .C(net300),
    .X(_1550_));
 sky130_fd_sc_hd__a221o_4 _3848_ (.A1(net2257),
    .A2(net239),
    .B1(net345),
    .B2(net241),
    .C1(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__inv_2 _3849_ (.A(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__xnor2_1 _3850_ (.A(_1549_),
    .B(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__mux4_1 _3851_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ),
    .A1(net39),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ),
    .S0(net364),
    .S1(net366),
    .X(_1554_));
 sky130_fd_sc_hd__a22o_1 _3852_ (.A1(net2217),
    .A2(net243),
    .B1(net344),
    .B2(_1345_),
    .X(_1555_));
 sky130_fd_sc_hd__a21oi_4 _3853_ (.A1(net2149),
    .A2(net304),
    .B1(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__mux2_2 _3854_ (.A0(_1300_),
    .A1(_1556_),
    .S(net363),
    .X(_1557_));
 sky130_fd_sc_hd__and3_1 _3855_ (.A(net2149),
    .B(_1356_),
    .C(_1360_),
    .X(_1558_));
 sky130_fd_sc_hd__a221o_4 _3856_ (.A1(net2294),
    .A2(net239),
    .B1(net344),
    .B2(net241),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__nand2_1 _3857_ (.A(_1539_),
    .B(_1542_),
    .Y(_1560_));
 sky130_fd_sc_hd__mux4_1 _3858_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ),
    .A1(net41),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ),
    .S0(net365),
    .S1(net367),
    .X(_1561_));
 sky130_fd_sc_hd__a22o_1 _3859_ (.A1(net2272),
    .A2(net242),
    .B1(net343),
    .B2(_1345_),
    .X(_1562_));
 sky130_fd_sc_hd__a21oi_2 _3860_ (.A1(net2198),
    .A2(net305),
    .B1(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_2 _3861_ (.A0(_1299_),
    .A1(_1563_),
    .S(net363),
    .X(_1564_));
 sky130_fd_sc_hd__and3_1 _3862_ (.A(net2198),
    .B(net332),
    .C(net301),
    .X(_1565_));
 sky130_fd_sc_hd__a221o_4 _3863_ (.A1(net2314),
    .A2(net239),
    .B1(net343),
    .B2(net240),
    .C1(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__or2_1 _3864_ (.A(_1564_),
    .B(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__o211a_1 _3865_ (.A1(_1557_),
    .A2(_1559_),
    .B1(_1560_),
    .C1(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__mux4_2 _3866_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ),
    .A1(net43),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ),
    .S0(net365),
    .S1(net367),
    .X(_1569_));
 sky130_fd_sc_hd__a22o_1 _3867_ (.A1(net2239),
    .A2(net242),
    .B1(net342),
    .B2(_1345_),
    .X(_1570_));
 sky130_fd_sc_hd__a21oi_4 _3868_ (.A1(net2023),
    .A2(net305),
    .B1(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__inv_2 _3869_ (.A(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__mux2_4 _3870_ (.A0(net2120),
    .A1(_1572_),
    .S(net362),
    .X(_1573_));
 sky130_fd_sc_hd__and3_1 _3871_ (.A(net2023),
    .B(net332),
    .C(net301),
    .X(_1574_));
 sky130_fd_sc_hd__a221o_4 _3872_ (.A1(net2296),
    .A2(net238),
    .B1(net342),
    .B2(net240),
    .C1(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__nand2b_1 _3873_ (.A_N(_1575_),
    .B(_1573_),
    .Y(_1576_));
 sky130_fd_sc_hd__xor2_1 _3874_ (.A(_1573_),
    .B(_1575_),
    .X(_1577_));
 sky130_fd_sc_hd__a21o_1 _3875_ (.A1(_1564_),
    .A2(_1566_),
    .B1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__mux4_2 _3876_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ),
    .A1(net40),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ),
    .S0(net364),
    .S1(net366),
    .X(_1579_));
 sky130_fd_sc_hd__and3_1 _3877_ (.A(net303),
    .B(net302),
    .C(net341),
    .X(_1580_));
 sky130_fd_sc_hd__a221o_4 _3878_ (.A1(net2012),
    .A2(net304),
    .B1(net243),
    .B2(net2275),
    .C1(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_2 _3879_ (.A0(net2199),
    .A1(_1581_),
    .S(net363),
    .X(_1582_));
 sky130_fd_sc_hd__and3_1 _3880_ (.A(net73),
    .B(net331),
    .C(net300),
    .X(_1583_));
 sky130_fd_sc_hd__a221o_4 _3881_ (.A1(net2340),
    .A2(net239),
    .B1(net341),
    .B2(net241),
    .C1(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__xor2_1 _3882_ (.A(_1582_),
    .B(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__a211oi_1 _3883_ (.A1(_1557_),
    .A2(_1559_),
    .B1(_1578_),
    .C1(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__and4bb_2 _3884_ (.A_N(_1544_),
    .B_N(_1553_),
    .C(_1568_),
    .D(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__mux4_2 _3885_ (.A0(net2353),
    .A1(net54),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ),
    .S0(net365),
    .S1(net367),
    .X(_1588_));
 sky130_fd_sc_hd__and3_1 _3886_ (.A(net303),
    .B(net302),
    .C(net340),
    .X(_1589_));
 sky130_fd_sc_hd__a221o_4 _3887_ (.A1(net2125),
    .A2(net305),
    .B1(net242),
    .B2(net2195),
    .C1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_2 _3888_ (.A0(net2310),
    .A1(_1590_),
    .S(net362),
    .X(_1591_));
 sky130_fd_sc_hd__inv_2 _3889_ (.A(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__and3_1 _3890_ (.A(net2125),
    .B(net332),
    .C(net301),
    .X(_1593_));
 sky130_fd_sc_hd__a221o_4 _3891_ (.A1(net2342),
    .A2(net238),
    .B1(net340),
    .B2(net240),
    .C1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__xor2_1 _3892_ (.A(_1591_),
    .B(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__mux4_2 _3893_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ),
    .A1(net52),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ),
    .S0(net365),
    .S1(net367),
    .X(_1596_));
 sky130_fd_sc_hd__a22o_1 _3894_ (.A1(net2181),
    .A2(net242),
    .B1(net339),
    .B2(_1345_),
    .X(_1597_));
 sky130_fd_sc_hd__a21oi_1 _3895_ (.A1(net85),
    .A2(net305),
    .B1(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__inv_2 _3896_ (.A(net2182),
    .Y(_1599_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(_1296_),
    .A1(_1598_),
    .S(net362),
    .X(_1600_));
 sky130_fd_sc_hd__mux2_1 _3898_ (.A0(net2173),
    .A1(_1599_),
    .S(net362),
    .X(_1601_));
 sky130_fd_sc_hd__and3_1 _3899_ (.A(net2186),
    .B(net332),
    .C(net301),
    .X(_1602_));
 sky130_fd_sc_hd__a221o_4 _3900_ (.A1(net2318),
    .A2(net238),
    .B1(net339),
    .B2(net240),
    .C1(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__a21o_1 _3901_ (.A1(_1600_),
    .A2(_1603_),
    .B1(_1595_),
    .X(_1604_));
 sky130_fd_sc_hd__mux4_2 _3902_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ),
    .A1(net49),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ),
    .S0(net365),
    .S1(net367),
    .X(_1605_));
 sky130_fd_sc_hd__and3_1 _3903_ (.A(net303),
    .B(net302),
    .C(net338),
    .X(_1606_));
 sky130_fd_sc_hd__a221o_2 _3904_ (.A1(net2024),
    .A2(net305),
    .B1(net242),
    .B2(net2300),
    .C1(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_2 _3905_ (.A0(net2155),
    .A1(_1607_),
    .S(net362),
    .X(_1608_));
 sky130_fd_sc_hd__inv_2 _3906_ (.A(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__and3_1 _3907_ (.A(net82),
    .B(net332),
    .C(net301),
    .X(_1610_));
 sky130_fd_sc_hd__a221o_4 _3908_ (.A1(net2320),
    .A2(net238),
    .B1(net338),
    .B2(net240),
    .C1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__xor2_1 _3909_ (.A(_1608_),
    .B(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__mux4_2 _3910_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ),
    .A1(net48),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ),
    .S0(net365),
    .S1(net367),
    .X(_1613_));
 sky130_fd_sc_hd__a22o_1 _3911_ (.A1(net549),
    .A2(net242),
    .B1(net337),
    .B2(_1345_),
    .X(_1614_));
 sky130_fd_sc_hd__a21oi_2 _3912_ (.A1(net537),
    .A2(net305),
    .B1(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__mux2_2 _3913_ (.A0(_1297_),
    .A1(_1615_),
    .S(net362),
    .X(_1616_));
 sky130_fd_sc_hd__and3_1 _3914_ (.A(net537),
    .B(net332),
    .C(net301),
    .X(_1617_));
 sky130_fd_sc_hd__a221o_4 _3915_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .A2(net238),
    .B1(net337),
    .B2(net240),
    .C1(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__a21o_1 _3916_ (.A1(_1616_),
    .A2(_1618_),
    .B1(_1612_),
    .X(_1619_));
 sky130_fd_sc_hd__nor2_1 _3917_ (.A(_1616_),
    .B(_1618_),
    .Y(_1620_));
 sky130_fd_sc_hd__or2_1 _3918_ (.A(_1600_),
    .B(_1603_),
    .X(_1621_));
 sky130_fd_sc_hd__mux4_2 _3919_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ),
    .A1(net50),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ),
    .S0(net365),
    .S1(net367),
    .X(_1622_));
 sky130_fd_sc_hd__and3_1 _3920_ (.A(net303),
    .B(net302),
    .C(net336),
    .X(_1623_));
 sky130_fd_sc_hd__a221o_4 _3921_ (.A1(net2143),
    .A2(net305),
    .B1(net242),
    .B2(net2250),
    .C1(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_2 _3922_ (.A0(net2289),
    .A1(_1624_),
    .S(net362),
    .X(_1625_));
 sky130_fd_sc_hd__and3_1 _3923_ (.A(net2143),
    .B(net332),
    .C(net301),
    .X(_1626_));
 sky130_fd_sc_hd__a221o_4 _3924_ (.A1(net2334),
    .A2(net238),
    .B1(net336),
    .B2(net240),
    .C1(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__and2b_1 _3925_ (.A_N(_1625_),
    .B(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__nand2b_1 _3926_ (.A_N(_1627_),
    .B(_1625_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_1621_),
    .B(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__or4_2 _3928_ (.A(_1619_),
    .B(_1620_),
    .C(_1628_),
    .D(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__mux4_2 _3929_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ),
    .A1(net55),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ),
    .S0(net365),
    .S1(net367),
    .X(_1632_));
 sky130_fd_sc_hd__and3_1 _3930_ (.A(net303),
    .B(net302),
    .C(net335),
    .X(_1633_));
 sky130_fd_sc_hd__a221o_4 _3931_ (.A1(net2163),
    .A2(net305),
    .B1(net242),
    .B2(net2196),
    .C1(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_2 _3932_ (.A0(net2297),
    .A1(_1634_),
    .S(net362),
    .X(_1635_));
 sky130_fd_sc_hd__and2_1 _3933_ (.A(net240),
    .B(net335),
    .X(_1636_));
 sky130_fd_sc_hd__a221oi_2 _3934_ (.A1(net88),
    .A2(_1361_),
    .B1(net238),
    .B2(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .C1(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__a221o_4 _3935_ (.A1(net2163),
    .A2(_1361_),
    .B1(net238),
    .B2(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .C1(_1636_),
    .X(_1638_));
 sky130_fd_sc_hd__or2_1 _3936_ (.A(_1635_),
    .B(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__nand2_1 _3937_ (.A(_1635_),
    .B(_1638_),
    .Y(_1640_));
 sky130_fd_sc_hd__and2_2 _3938_ (.A(_1639_),
    .B(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__mux4_2 _3939_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ),
    .A1(net47),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ),
    .S0(net365),
    .S1(net367),
    .X(_1642_));
 sky130_fd_sc_hd__a22o_1 _3940_ (.A1(net2279),
    .A2(net243),
    .B1(_1642_),
    .B2(_1345_),
    .X(_1643_));
 sky130_fd_sc_hd__a21oi_4 _3941_ (.A1(net2103),
    .A2(net304),
    .B1(net2280),
    .Y(_1644_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(net2302),
    .B(net2240),
    .Y(_1645_));
 sky130_fd_sc_hd__o21ai_4 _3943_ (.A1(net2302),
    .A2(_1644_),
    .B1(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__and3_1 _3944_ (.A(net80),
    .B(net332),
    .C(net301),
    .X(_1647_));
 sky130_fd_sc_hd__a221o_4 _3945_ (.A1(net2330),
    .A2(net238),
    .B1(net334),
    .B2(net240),
    .C1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__inv_2 _3946_ (.A(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__xnor2_1 _3947_ (.A(_1646_),
    .B(_1648_),
    .Y(_1650_));
 sky130_fd_sc_hd__mux4_2 _3948_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ),
    .A1(net51),
    .A2(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ),
    .S0(net365),
    .S1(net367),
    .X(_1651_));
 sky130_fd_sc_hd__and3_1 _3949_ (.A(net303),
    .B(net302),
    .C(net333),
    .X(_1652_));
 sky130_fd_sc_hd__a221o_1 _3950_ (.A1(net1704),
    .A2(net305),
    .B1(net242),
    .B2(net2207),
    .C1(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_2 _3951_ (.A0(net2183),
    .A1(_1653_),
    .S(net362),
    .X(_1654_));
 sky130_fd_sc_hd__and3_1 _3952_ (.A(net84),
    .B(net332),
    .C(net301),
    .X(_1655_));
 sky130_fd_sc_hd__a221o_4 _3953_ (.A1(net2341),
    .A2(net238),
    .B1(net333),
    .B2(net240),
    .C1(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__xnor2_1 _3954_ (.A(_1654_),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__inv_2 _3955_ (.A(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_1 _3956_ (.A(_1650_),
    .B(_1657_),
    .Y(_1659_));
 sky130_fd_sc_hd__nor4_4 _3957_ (.A(_1604_),
    .B(_1631_),
    .C(_1641_),
    .D(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand4_4 _3958_ (.A(_1419_),
    .B(_1518_),
    .C(_1587_),
    .D(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__o211ai_2 _3959_ (.A1(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .A2(_1474_),
    .B1(_1475_),
    .C1(_1478_),
    .Y(_1662_));
 sky130_fd_sc_hd__a21o_1 _3960_ (.A1(net204),
    .A2(_1662_),
    .B1(_1443_),
    .X(_1663_));
 sky130_fd_sc_hd__or2_1 _3961_ (.A(net204),
    .B(_1662_),
    .X(_1664_));
 sky130_fd_sc_hd__inv_2 _3962_ (.A(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__nor2_1 _3963_ (.A(net201),
    .B(_1469_),
    .Y(_1666_));
 sky130_fd_sc_hd__a311o_1 _3964_ (.A1(_1470_),
    .A2(_1663_),
    .A3(_1664_),
    .B1(_1666_),
    .C1(_1452_),
    .X(_1667_));
 sky130_fd_sc_hd__nor2_1 _3965_ (.A(net217),
    .B(_1427_),
    .Y(_1668_));
 sky130_fd_sc_hd__a211o_1 _3966_ (.A1(_1438_),
    .A2(_1667_),
    .B1(_1668_),
    .C1(_1460_),
    .X(_1669_));
 sky130_fd_sc_hd__and3b_1 _3967_ (.A_N(_1488_),
    .B(_1497_),
    .C(_1486_),
    .X(_1670_));
 sky130_fd_sc_hd__a221o_1 _3968_ (.A1(_1493_),
    .A2(_1496_),
    .B1(_1500_),
    .B2(_1669_),
    .C1(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__a21o_1 _3969_ (.A1(_1354_),
    .A2(_1372_),
    .B1(_1391_),
    .X(_1672_));
 sky130_fd_sc_hd__o211a_1 _3970_ (.A1(_1399_),
    .A2(_1408_),
    .B1(_1418_),
    .C1(_1400_),
    .X(_1673_));
 sky130_fd_sc_hd__and2b_1 _3971_ (.A_N(_1417_),
    .B(_1415_),
    .X(_1674_));
 sky130_fd_sc_hd__o31a_1 _3972_ (.A1(_1383_),
    .A2(_1673_),
    .A3(_1674_),
    .B1(_1382_),
    .X(_1675_));
 sky130_fd_sc_hd__a211o_1 _3973_ (.A1(_1419_),
    .A2(_1671_),
    .B1(_1672_),
    .C1(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__and3b_1 _3974_ (.A_N(_1506_),
    .B(_1514_),
    .C(_1504_),
    .X(_1677_));
 sky130_fd_sc_hd__a211o_1 _3975_ (.A1(_1517_),
    .A2(_1676_),
    .B1(_1677_),
    .C1(_1515_),
    .X(_1678_));
 sky130_fd_sc_hd__a21oi_1 _3976_ (.A1(_1530_),
    .A2(_1533_),
    .B1(_1524_),
    .Y(_1679_));
 sky130_fd_sc_hd__a21o_1 _3977_ (.A1(_1522_),
    .A2(_1679_),
    .B1(_1534_),
    .X(_1680_));
 sky130_fd_sc_hd__o2bb2a_1 _3978_ (.A1_N(_1549_),
    .A2_N(_1552_),
    .B1(_1557_),
    .B2(_1559_),
    .X(_1681_));
 sky130_fd_sc_hd__a211o_1 _3979_ (.A1(_1557_),
    .A2(_1559_),
    .B1(_1585_),
    .C1(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__nand2b_1 _3980_ (.A_N(_1584_),
    .B(_1582_),
    .Y(_1683_));
 sky130_fd_sc_hd__a31o_1 _3981_ (.A1(_1567_),
    .A2(_1682_),
    .A3(_1683_),
    .B1(_1578_),
    .X(_1684_));
 sky130_fd_sc_hd__a31oi_2 _3982_ (.A1(_1560_),
    .A2(_1576_),
    .A3(_1684_),
    .B1(_1544_),
    .Y(_1685_));
 sky130_fd_sc_hd__a211o_1 _3983_ (.A1(_1587_),
    .A2(_1678_),
    .B1(_1680_),
    .C1(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__a21oi_1 _3984_ (.A1(_1646_),
    .A2(_1649_),
    .B1(_1620_),
    .Y(_1687_));
 sky130_fd_sc_hd__o221a_1 _3985_ (.A1(_1609_),
    .A2(_1611_),
    .B1(_1619_),
    .B2(_1687_),
    .C1(_1629_),
    .X(_1688_));
 sky130_fd_sc_hd__nand2b_1 _3986_ (.A_N(_1656_),
    .B(_1654_),
    .Y(_1689_));
 sky130_fd_sc_hd__o311a_1 _3987_ (.A1(_1628_),
    .A2(_1658_),
    .A3(_1688_),
    .B1(_1689_),
    .C1(_1621_),
    .X(_1690_));
 sky130_fd_sc_hd__o22a_1 _3988_ (.A1(_1592_),
    .A2(_1594_),
    .B1(_1604_),
    .B2(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__nor2_1 _3989_ (.A(_1641_),
    .B(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__a221o_1 _3990_ (.A1(_1635_),
    .A2(net190),
    .B1(_1660_),
    .B2(_1686_),
    .C1(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__and3_1 _3991_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(_1661_),
    .C(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .Y(_1695_));
 sky130_fd_sc_hd__a21oi_1 _3993_ (.A1(_1661_),
    .A2(_1693_),
    .B1(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .Y(_1696_));
 sky130_fd_sc_hd__or4_1 _3994_ (.A(net2238),
    .B(_1694_),
    .C(_1695_),
    .D(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__nand2b_2 _3995_ (.A_N(net2292),
    .B(net2251),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(net2252),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2b_4 _3997_ (.A_N(net2251),
    .B(net2292),
    .Y(_1700_));
 sky130_fd_sc_hd__or2_2 _3998_ (.A(net2252),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(_1701_));
 sky130_fd_sc_hd__a221o_1 _3999_ (.A1(_1698_),
    .A2(net2253),
    .B1(_1700_),
    .B2(_1701_),
    .C1(net2208),
    .X(_1702_));
 sky130_fd_sc_hd__or3b_4 _4000_ (.A(net2252),
    .B(net2208),
    .C_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(_1703_));
 sky130_fd_sc_hd__o21a_1 _4001_ (.A1(_1698_),
    .A2(_1703_),
    .B1(_1702_),
    .X(_1704_));
 sky130_fd_sc_hd__or3_1 _4002_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .B(_1698_),
    .C(_1699_),
    .X(_1705_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(_1704_),
    .A1(_1705_),
    .S(_1661_),
    .X(_1706_));
 sky130_fd_sc_hd__a21bo_1 _4004_ (.A1(_1697_),
    .A2(_1706_),
    .B1_N(net2130),
    .X(_1707_));
 sky130_fd_sc_hd__and2_1 _4005_ (.A(_1301_),
    .B(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__mux2_1 _4006_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .S(net428),
    .X(_1709_));
 sky130_fd_sc_hd__xnor2_1 _4007_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .B(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__mux2_1 _4008_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .S(net428),
    .X(_1711_));
 sky130_fd_sc_hd__nand2_1 _4009_ (.A(net2173),
    .B(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__or2_1 _4010_ (.A(net2173),
    .B(_1711_),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_1 _4011_ (.A(net2174),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__mux2_1 _4012_ (.A0(net2218),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .S(net428),
    .X(_1715_));
 sky130_fd_sc_hd__nand2_1 _4013_ (.A(net2183),
    .B(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__or2_1 _4014_ (.A(net2183),
    .B(net2219),
    .X(_1717_));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(net2184),
    .B(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__mux2_1 _4016_ (.A0(net2159),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .S(net428),
    .X(_1719_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .B(net2160),
    .Y(_1720_));
 sky130_fd_sc_hd__or2_1 _4018_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .B(net2160),
    .X(_1721_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(net2161),
    .B(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__mux2_1 _4020_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ),
    .A1(net2351),
    .S(net428),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(net2155),
    .B(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__or2_1 _4022_ (.A(net2155),
    .B(_1723_),
    .X(_1725_));
 sky130_fd_sc_hd__nand2_1 _4023_ (.A(net2156),
    .B(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .S(net428),
    .X(_1727_));
 sky130_fd_sc_hd__nand2_1 _4025_ (.A(net2113),
    .B(_1727_),
    .Y(_1728_));
 sky130_fd_sc_hd__or2_1 _4026_ (.A(net2113),
    .B(_1727_),
    .X(_1729_));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(net2114),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(net2203),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .S(net428),
    .X(_1731_));
 sky130_fd_sc_hd__xnor2_1 _4029_ (.A(net2240),
    .B(net2204),
    .Y(_1732_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .S(net428),
    .X(_1733_));
 sky130_fd_sc_hd__and2_1 _4031_ (.A(net2177),
    .B(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__nor2_1 _4032_ (.A(net2177),
    .B(_1733_),
    .Y(_1735_));
 sky130_fd_sc_hd__or2_1 _4033_ (.A(_1734_),
    .B(net2178),
    .X(_1736_));
 sky130_fd_sc_hd__mux2_1 _4034_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .S(net428),
    .X(_1737_));
 sky130_fd_sc_hd__and2_1 _4035_ (.A(net2151),
    .B(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__nor2_1 _4036_ (.A(net2151),
    .B(_1737_),
    .Y(_1739_));
 sky130_fd_sc_hd__or2_1 _4037_ (.A(_1738_),
    .B(net2152),
    .X(_1740_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .S(net428),
    .X(_1741_));
 sky130_fd_sc_hd__and2_1 _4039_ (.A(net2077),
    .B(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__nor2_1 _4040_ (.A(net2077),
    .B(_1741_),
    .Y(_1743_));
 sky130_fd_sc_hd__or2_1 _4041_ (.A(_1742_),
    .B(net2078),
    .X(_1744_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .S(net428),
    .X(_1745_));
 sky130_fd_sc_hd__and2_1 _4043_ (.A(net2120),
    .B(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__nor2_1 _4044_ (.A(net2120),
    .B(_1745_),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _4045_ (.A(_1746_),
    .B(net2121),
    .X(_1748_));
 sky130_fd_sc_hd__mux2_1 _4046_ (.A0(net2319),
    .A1(net2314),
    .S(net428),
    .X(_1749_));
 sky130_fd_sc_hd__and2_2 _4047_ (.A(net2306),
    .B(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__nor2_1 _4048_ (.A(net2306),
    .B(_1749_),
    .Y(_1751_));
 sky130_fd_sc_hd__or2_1 _4049_ (.A(net2307),
    .B(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .S(net427),
    .X(_1753_));
 sky130_fd_sc_hd__and2_1 _4051_ (.A(net2199),
    .B(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__nor2_1 _4052_ (.A(net2199),
    .B(_1753_),
    .Y(_1755_));
 sky130_fd_sc_hd__or2_1 _4053_ (.A(_1754_),
    .B(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .S(net427),
    .X(_1757_));
 sky130_fd_sc_hd__and2_1 _4055_ (.A(net2317),
    .B(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__nor2_1 _4056_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .B(_1757_),
    .Y(_1759_));
 sky130_fd_sc_hd__or2_1 _4057_ (.A(_1758_),
    .B(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .S(net428),
    .X(_1761_));
 sky130_fd_sc_hd__and2_1 _4059_ (.A(net2134),
    .B(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__nor2_1 _4060_ (.A(net2134),
    .B(_1761_),
    .Y(_1763_));
 sky130_fd_sc_hd__or2_1 _4061_ (.A(net2135),
    .B(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(net2242),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .S(net427),
    .X(_1765_));
 sky130_fd_sc_hd__and2_1 _4063_ (.A(net2088),
    .B(net2243),
    .X(_1766_));
 sky130_fd_sc_hd__nor2_1 _4064_ (.A(net2088),
    .B(_1765_),
    .Y(_1767_));
 sky130_fd_sc_hd__or2_1 _4065_ (.A(_1766_),
    .B(net2089),
    .X(_1768_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .S(net427),
    .X(_1769_));
 sky130_fd_sc_hd__and2_1 _4067_ (.A(net2224),
    .B(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__nor2_1 _4068_ (.A(net2224),
    .B(_1769_),
    .Y(_1771_));
 sky130_fd_sc_hd__or2_1 _4069_ (.A(net2225),
    .B(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__mux2_1 _4070_ (.A0(net2270),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .S(net427),
    .X(_1773_));
 sky130_fd_sc_hd__and2_1 _4071_ (.A(net2171),
    .B(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__nor2_1 _4072_ (.A(net2171),
    .B(_1773_),
    .Y(_1775_));
 sky130_fd_sc_hd__or2_1 _4073_ (.A(_1774_),
    .B(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .S(net427),
    .X(_1777_));
 sky130_fd_sc_hd__and2_1 _4075_ (.A(net2098),
    .B(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__nor2_1 _4076_ (.A(net2098),
    .B(_1777_),
    .Y(_1779_));
 sky130_fd_sc_hd__or2_1 _4077_ (.A(_1778_),
    .B(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ),
    .S(net427),
    .X(_1781_));
 sky130_fd_sc_hd__and2_1 _4079_ (.A(net2205),
    .B(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__nor2_1 _4080_ (.A(net2205),
    .B(_1781_),
    .Y(_1783_));
 sky130_fd_sc_hd__or2_1 _4081_ (.A(net2206),
    .B(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__mux2_1 _4082_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .S(net427),
    .X(_1785_));
 sky130_fd_sc_hd__and2_1 _4083_ (.A(net2211),
    .B(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__nor2_1 _4084_ (.A(net2211),
    .B(_1785_),
    .Y(_1787_));
 sky130_fd_sc_hd__or2_1 _4085_ (.A(_1786_),
    .B(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__mux2_2 _4086_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .S(net427),
    .X(_1789_));
 sky130_fd_sc_hd__and2_1 _4087_ (.A(net2215),
    .B(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__nor2_1 _4088_ (.A(net2215),
    .B(_1789_),
    .Y(_1791_));
 sky130_fd_sc_hd__or2_1 _4089_ (.A(_1790_),
    .B(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(net2230),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .S(net427),
    .X(_1793_));
 sky130_fd_sc_hd__and2_1 _4091_ (.A(net2138),
    .B(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__nor2_1 _4092_ (.A(net2138),
    .B(_1793_),
    .Y(_1795_));
 sky130_fd_sc_hd__or2_1 _4093_ (.A(_1794_),
    .B(net2139),
    .X(_1796_));
 sky130_fd_sc_hd__mux2_1 _4094_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .S(net427),
    .X(_1797_));
 sky130_fd_sc_hd__and2_1 _4095_ (.A(net2188),
    .B(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__nor2_1 _4096_ (.A(net2188),
    .B(_1797_),
    .Y(_1799_));
 sky130_fd_sc_hd__or2_1 _4097_ (.A(_1798_),
    .B(net2189),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_2 _4098_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .S(net427),
    .X(_1801_));
 sky130_fd_sc_hd__and2_1 _4099_ (.A(net2235),
    .B(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__nor2_1 _4100_ (.A(net2235),
    .B(_1801_),
    .Y(_1803_));
 sky130_fd_sc_hd__or2_1 _4101_ (.A(_1802_),
    .B(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .S(net427),
    .X(_1805_));
 sky130_fd_sc_hd__and2_1 _4103_ (.A(net2067),
    .B(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__nor2_1 _4104_ (.A(net2067),
    .B(_1805_),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_1 _4105_ (.A(_1806_),
    .B(net2068),
    .X(_1808_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .S(net427),
    .X(_1809_));
 sky130_fd_sc_hd__and2_1 _4107_ (.A(net2273),
    .B(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__nor2_1 _4108_ (.A(net2273),
    .B(_1809_),
    .Y(_1811_));
 sky130_fd_sc_hd__or2_1 _4109_ (.A(net2274),
    .B(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(net2276),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .S(net427),
    .X(_1813_));
 sky130_fd_sc_hd__and2_1 _4111_ (.A(net2107),
    .B(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__nor2_1 _4112_ (.A(net2107),
    .B(_1813_),
    .Y(_1815_));
 sky130_fd_sc_hd__or2_1 _4113_ (.A(_1814_),
    .B(net2108),
    .X(_1816_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .S(net428),
    .X(_1817_));
 sky130_fd_sc_hd__and2_1 _4115_ (.A(net2226),
    .B(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__and3_1 _4116_ (.A(net826),
    .B(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .C(net2282),
    .X(_1819_));
 sky130_fd_sc_hd__a21oi_1 _4117_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .A2(net427),
    .B1(net826),
    .Y(_1820_));
 sky130_fd_sc_hd__or2_1 _4118_ (.A(_1819_),
    .B(net827),
    .X(_1821_));
 sky130_fd_sc_hd__nand3_1 _4119_ (.A(net773),
    .B(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .C(net2282),
    .Y(_1822_));
 sky130_fd_sc_hd__nor2_1 _4120_ (.A(net828),
    .B(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__nor2_1 _4121_ (.A(net2226),
    .B(_1817_),
    .Y(_1824_));
 sky130_fd_sc_hd__or2_1 _4122_ (.A(_1818_),
    .B(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__o21ba_1 _4123_ (.A1(net2283),
    .A2(_1823_),
    .B1_N(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__nor2_1 _4124_ (.A(_1818_),
    .B(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__o21ba_1 _4125_ (.A1(_1818_),
    .A2(_1826_),
    .B1_N(_1816_),
    .X(_1828_));
 sky130_fd_sc_hd__or2_1 _4126_ (.A(_1814_),
    .B(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__o21ba_1 _4127_ (.A1(_1814_),
    .A2(_1828_),
    .B1_N(_1812_),
    .X(_1830_));
 sky130_fd_sc_hd__or2_1 _4128_ (.A(_1810_),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__o21ba_1 _4129_ (.A1(_1810_),
    .A2(_1830_),
    .B1_N(_1808_),
    .X(_1832_));
 sky130_fd_sc_hd__or2_1 _4130_ (.A(_1806_),
    .B(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__o21ba_1 _4131_ (.A1(_1806_),
    .A2(_1832_),
    .B1_N(_1804_),
    .X(_1834_));
 sky130_fd_sc_hd__or2_1 _4132_ (.A(_1802_),
    .B(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__o21ba_1 _4133_ (.A1(_1802_),
    .A2(_1834_),
    .B1_N(_1800_),
    .X(_1836_));
 sky130_fd_sc_hd__nor2_1 _4134_ (.A(_1798_),
    .B(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__o21ba_1 _4135_ (.A1(_1798_),
    .A2(_1836_),
    .B1_N(_1796_),
    .X(_1838_));
 sky130_fd_sc_hd__or2_1 _4136_ (.A(_1794_),
    .B(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__o21ba_1 _4137_ (.A1(_1794_),
    .A2(_1838_),
    .B1_N(_1792_),
    .X(_1840_));
 sky130_fd_sc_hd__or2_1 _4138_ (.A(_1790_),
    .B(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__o21ba_1 _4139_ (.A1(_1790_),
    .A2(_1840_),
    .B1_N(_1788_),
    .X(_1842_));
 sky130_fd_sc_hd__nor2_1 _4140_ (.A(net2212),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__o21ba_1 _4141_ (.A1(_1786_),
    .A2(_1842_),
    .B1_N(_1784_),
    .X(_1844_));
 sky130_fd_sc_hd__or2_1 _4142_ (.A(_1782_),
    .B(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__o21ba_1 _4143_ (.A1(_1782_),
    .A2(_1844_),
    .B1_N(_1780_),
    .X(_1846_));
 sky130_fd_sc_hd__or2_1 _4144_ (.A(_1778_),
    .B(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__o21ba_1 _4145_ (.A1(_1778_),
    .A2(_1846_),
    .B1_N(_1776_),
    .X(_1848_));
 sky130_fd_sc_hd__nor2_1 _4146_ (.A(_1774_),
    .B(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__o21ba_1 _4147_ (.A1(_1774_),
    .A2(_1848_),
    .B1_N(_1772_),
    .X(_1850_));
 sky130_fd_sc_hd__or2_1 _4148_ (.A(_1770_),
    .B(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__o21ba_1 _4149_ (.A1(_1770_),
    .A2(_1850_),
    .B1_N(_1768_),
    .X(_1852_));
 sky130_fd_sc_hd__or2_1 _4150_ (.A(_1766_),
    .B(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__o21ba_1 _4151_ (.A1(_1766_),
    .A2(_1852_),
    .B1_N(_1764_),
    .X(_1854_));
 sky130_fd_sc_hd__or2_1 _4152_ (.A(net2135),
    .B(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o21ba_1 _4153_ (.A1(_1762_),
    .A2(_1854_),
    .B1_N(_1760_),
    .X(_1856_));
 sky130_fd_sc_hd__or2_1 _4154_ (.A(_1758_),
    .B(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__o21ba_1 _4155_ (.A1(_1758_),
    .A2(_1856_),
    .B1_N(_1756_),
    .X(_1858_));
 sky130_fd_sc_hd__or2_1 _4156_ (.A(_1754_),
    .B(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__o21ba_2 _4157_ (.A1(_1754_),
    .A2(_1858_),
    .B1_N(_1752_),
    .X(_1860_));
 sky130_fd_sc_hd__nor2_1 _4158_ (.A(_1750_),
    .B(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__o21ba_1 _4159_ (.A1(_1750_),
    .A2(_1860_),
    .B1_N(_1748_),
    .X(_1862_));
 sky130_fd_sc_hd__or2_1 _4160_ (.A(_1746_),
    .B(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__o21ba_1 _4161_ (.A1(_1746_),
    .A2(_1862_),
    .B1_N(_1744_),
    .X(_1864_));
 sky130_fd_sc_hd__or2_1 _4162_ (.A(_1742_),
    .B(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__o21ba_1 _4163_ (.A1(_1742_),
    .A2(_1864_),
    .B1_N(_1740_),
    .X(_1866_));
 sky130_fd_sc_hd__nor2_1 _4164_ (.A(_1738_),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__o21ba_1 _4165_ (.A1(_1738_),
    .A2(_1866_),
    .B1_N(_1736_),
    .X(_1868_));
 sky130_fd_sc_hd__or2_1 _4166_ (.A(_1734_),
    .B(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__o21ba_1 _4167_ (.A1(_1734_),
    .A2(_1868_),
    .B1_N(_1732_),
    .X(_1870_));
 sky130_fd_sc_hd__a21oi_2 _4168_ (.A1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .A2(_1731_),
    .B1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__o21a_1 _4169_ (.A1(_1730_),
    .A2(_1871_),
    .B1(net2114),
    .X(_1872_));
 sky130_fd_sc_hd__o21a_1 _4170_ (.A1(_1726_),
    .A2(_1872_),
    .B1(net2156),
    .X(_1873_));
 sky130_fd_sc_hd__o21a_1 _4171_ (.A1(_1722_),
    .A2(_1873_),
    .B1(net2161),
    .X(_1874_));
 sky130_fd_sc_hd__o21a_1 _4172_ (.A1(_1718_),
    .A2(_1874_),
    .B1(net2184),
    .X(_1875_));
 sky130_fd_sc_hd__o21ai_1 _4173_ (.A1(_1714_),
    .A2(_1875_),
    .B1(net2174),
    .Y(_1876_));
 sky130_fd_sc_hd__and2b_1 _4174_ (.A_N(_1710_),
    .B(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__a21oi_1 _4175_ (.A1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .A2(_1709_),
    .B1(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__xnor2_2 _4176_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .B(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(net2227),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .S(net428),
    .X(_1880_));
 sky130_fd_sc_hd__xor2_1 _4178_ (.A(_1879_),
    .B(net2228),
    .X(_1881_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(net2229),
    .A1(net2041),
    .S(net184),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(net2150),
    .A1(_1882_),
    .S(net247),
    .X(_1274_));
 sky130_fd_sc_hd__xnor2_1 _4181_ (.A(_1710_),
    .B(net2175),
    .Y(_1883_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(net2176),
    .A1(net2061),
    .S(net184),
    .X(_1884_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(net2064),
    .A1(_1884_),
    .S(net245),
    .X(_1273_));
 sky130_fd_sc_hd__xnor2_1 _4184_ (.A(_1714_),
    .B(_1875_),
    .Y(_1885_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(_1886_),
    .A1(net2051),
    .S(net184),
    .X(_1887_));
 sky130_fd_sc_hd__mux2_1 _4187_ (.A0(net1696),
    .A1(_1887_),
    .S(net244),
    .X(_1272_));
 sky130_fd_sc_hd__xnor2_1 _4188_ (.A(_1718_),
    .B(_1874_),
    .Y(_1888_));
 sky130_fd_sc_hd__inv_2 _4189_ (.A(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(_1889_),
    .A1(net2025),
    .S(net184),
    .X(_1890_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(net2005),
    .A1(_1890_),
    .S(net244),
    .X(_1271_));
 sky130_fd_sc_hd__xnor2_2 _4192_ (.A(net2162),
    .B(_1873_),
    .Y(_1891_));
 sky130_fd_sc_hd__inv_2 _4193_ (.A(_1891_),
    .Y(_1892_));
 sky130_fd_sc_hd__mux2_2 _4194_ (.A0(_1892_),
    .A1(net2066),
    .S(net184),
    .X(_1893_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net2194),
    .A1(_1893_),
    .S(net244),
    .X(_1270_));
 sky130_fd_sc_hd__xnor2_1 _4196_ (.A(net2157),
    .B(_1872_),
    .Y(_1894_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(_1895_),
    .A1(net1955),
    .S(net184),
    .X(_1896_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net2003),
    .A1(_1896_),
    .S(net247),
    .X(_1269_));
 sky130_fd_sc_hd__xnor2_1 _4200_ (.A(net2115),
    .B(_1871_),
    .Y(_1897_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(net2116),
    .Y(_1898_));
 sky130_fd_sc_hd__mux2_2 _4202_ (.A0(_1898_),
    .A1(net2036),
    .S(net184),
    .X(_1899_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(net834),
    .A1(_1899_),
    .S(net246),
    .X(_1268_));
 sky130_fd_sc_hd__xnor2_1 _4204_ (.A(_1732_),
    .B(_1869_),
    .Y(_1900_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(_1900_),
    .A1(net2047),
    .S(net2209),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(net2071),
    .A1(_1901_),
    .S(net246),
    .X(_1267_));
 sky130_fd_sc_hd__xnor2_1 _4207_ (.A(net2179),
    .B(_1867_),
    .Y(_1902_));
 sky130_fd_sc_hd__inv_2 _4208_ (.A(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(_1903_),
    .A1(net2073),
    .S(net184),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(net1711),
    .A1(_1904_),
    .S(net244),
    .X(_1266_));
 sky130_fd_sc_hd__xnor2_1 _4211_ (.A(net2153),
    .B(_1865_),
    .Y(_1905_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(_1905_),
    .A1(net2060),
    .S(net184),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(net2165),
    .A1(_1906_),
    .S(net244),
    .X(_1265_));
 sky130_fd_sc_hd__xnor2_1 _4214_ (.A(net2079),
    .B(_1863_),
    .Y(_1907_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(_1907_),
    .A1(net2033),
    .S(net184),
    .X(_1908_));
 sky130_fd_sc_hd__mux2_1 _4216_ (.A0(net2142),
    .A1(net2081),
    .S(net246),
    .X(_1264_));
 sky130_fd_sc_hd__xnor2_1 _4217_ (.A(net2122),
    .B(_1861_),
    .Y(_1909_));
 sky130_fd_sc_hd__inv_2 _4218_ (.A(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(_1910_),
    .A1(net2007),
    .S(net184),
    .X(_1911_));
 sky130_fd_sc_hd__inv_2 _4220_ (.A(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(net786),
    .A1(net2124),
    .S(net246),
    .X(_1263_));
 sky130_fd_sc_hd__xnor2_1 _4222_ (.A(_1752_),
    .B(_1859_),
    .Y(_1913_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(_1913_),
    .A1(net2049),
    .S(net184),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(net1973),
    .A1(net2050),
    .S(net250),
    .X(_1262_));
 sky130_fd_sc_hd__xnor2_1 _4225_ (.A(_1756_),
    .B(_1857_),
    .Y(_1915_));
 sky130_fd_sc_hd__mux2_2 _4226_ (.A0(_1915_),
    .A1(net889),
    .S(net183),
    .X(_1916_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(net1948),
    .A1(_1916_),
    .S(net252),
    .X(_1261_));
 sky130_fd_sc_hd__xnor2_1 _4228_ (.A(_1760_),
    .B(net2136),
    .Y(_1917_));
 sky130_fd_sc_hd__mux2_1 _4229_ (.A0(net2137),
    .A1(net2034),
    .S(net184),
    .X(_1918_));
 sky130_fd_sc_hd__mux2_1 _4230_ (.A0(net1034),
    .A1(_1918_),
    .S(net249),
    .X(_1260_));
 sky130_fd_sc_hd__xnor2_1 _4231_ (.A(_1764_),
    .B(_1853_),
    .Y(_1919_));
 sky130_fd_sc_hd__mux2_2 _4232_ (.A0(_1919_),
    .A1(net2062),
    .S(net183),
    .X(_1920_));
 sky130_fd_sc_hd__mux2_1 _4233_ (.A0(net2072),
    .A1(_1920_),
    .S(net250),
    .X(_1259_));
 sky130_fd_sc_hd__xnor2_1 _4234_ (.A(net2090),
    .B(_1851_),
    .Y(_1921_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(_1921_),
    .A1(net2083),
    .S(net183),
    .X(_1922_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(net2013),
    .A1(_1922_),
    .S(net251),
    .X(_1258_));
 sky130_fd_sc_hd__xnor2_1 _4237_ (.A(_1772_),
    .B(_1849_),
    .Y(_1923_));
 sky130_fd_sc_hd__inv_2 _4238_ (.A(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__mux2_2 _4239_ (.A0(_1924_),
    .A1(net2009),
    .S(net183),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(net2014),
    .A1(_1925_),
    .S(net252),
    .X(_1257_));
 sky130_fd_sc_hd__xnor2_1 _4241_ (.A(_1776_),
    .B(_1847_),
    .Y(_1926_));
 sky130_fd_sc_hd__mux2_2 _4242_ (.A0(_1926_),
    .A1(net2027),
    .S(net183),
    .X(_1927_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(net1811),
    .A1(net2028),
    .S(net250),
    .X(_1256_));
 sky130_fd_sc_hd__xnor2_1 _4244_ (.A(_1780_),
    .B(_1845_),
    .Y(_1928_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(_1928_),
    .A1(net1741),
    .S(net183),
    .X(_1929_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(net627),
    .A1(_1929_),
    .S(net253),
    .X(_1255_));
 sky130_fd_sc_hd__xnor2_1 _4247_ (.A(_1784_),
    .B(net2213),
    .Y(_1930_));
 sky130_fd_sc_hd__inv_2 _4248_ (.A(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__mux2_2 _4249_ (.A0(_1931_),
    .A1(net2065),
    .S(net183),
    .X(_1932_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(net2004),
    .A1(_1932_),
    .S(net251),
    .X(_1254_));
 sky130_fd_sc_hd__xnor2_2 _4251_ (.A(_1788_),
    .B(_1841_),
    .Y(_1933_));
 sky130_fd_sc_hd__mux2_4 _4252_ (.A0(_1933_),
    .A1(net2043),
    .S(net184),
    .X(_1934_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(net1966),
    .A1(_1934_),
    .S(net248),
    .X(_1253_));
 sky130_fd_sc_hd__xnor2_2 _4254_ (.A(_1792_),
    .B(_1839_),
    .Y(_1935_));
 sky130_fd_sc_hd__mux2_2 _4255_ (.A0(_1935_),
    .A1(net2016),
    .S(net183),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(net795),
    .A1(_1936_),
    .S(net252),
    .X(_1252_));
 sky130_fd_sc_hd__xnor2_1 _4257_ (.A(net2140),
    .B(_1837_),
    .Y(_1937_));
 sky130_fd_sc_hd__inv_2 _4258_ (.A(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__mux2_2 _4259_ (.A0(_1938_),
    .A1(net2017),
    .S(net183),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(net1758),
    .A1(_1939_),
    .S(net249),
    .X(_1251_));
 sky130_fd_sc_hd__xnor2_1 _4261_ (.A(net2190),
    .B(_1835_),
    .Y(_1940_));
 sky130_fd_sc_hd__mux2_2 _4262_ (.A0(_1940_),
    .A1(net949),
    .S(net183),
    .X(_1941_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net768),
    .A1(_1941_),
    .S(net249),
    .X(_1250_));
 sky130_fd_sc_hd__xnor2_1 _4264_ (.A(_1804_),
    .B(_1833_),
    .Y(_1942_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(_1942_),
    .A1(net1998),
    .S(net183),
    .X(_1943_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(net577),
    .A1(_1943_),
    .S(net250),
    .X(_1249_));
 sky130_fd_sc_hd__xnor2_1 _4267_ (.A(net2069),
    .B(_1831_),
    .Y(_1944_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(_1944_),
    .A1(net2008),
    .S(net183),
    .X(_1945_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net2075),
    .A1(_1945_),
    .S(net251),
    .X(_1248_));
 sky130_fd_sc_hd__xnor2_1 _4270_ (.A(_1812_),
    .B(_1829_),
    .Y(_1946_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(_1946_),
    .A1(net2015),
    .S(net183),
    .X(_1947_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(net2147),
    .A1(_1947_),
    .S(net251),
    .X(_1247_));
 sky130_fd_sc_hd__xnor2_1 _4273_ (.A(net2109),
    .B(_1827_),
    .Y(_1948_));
 sky130_fd_sc_hd__inv_2 _4274_ (.A(_1948_),
    .Y(_1949_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(_1949_),
    .A1(net2040),
    .S(net183),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(net1324),
    .A1(_1950_),
    .S(net252),
    .X(_1246_));
 sky130_fd_sc_hd__or3b_1 _4277_ (.A(net2283),
    .B(_1823_),
    .C_N(_1825_),
    .X(_1951_));
 sky130_fd_sc_hd__nand2b_1 _4278_ (.A_N(_1826_),
    .B(net2284),
    .Y(_1952_));
 sky130_fd_sc_hd__inv_2 _4279_ (.A(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(_1953_),
    .A1(net2082),
    .S(net183),
    .X(_1954_));
 sky130_fd_sc_hd__nor2_1 _4281_ (.A(net264),
    .B(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__o21ba_1 _4282_ (.A1(net978),
    .A2(net250),
    .B1_N(_1955_),
    .X(_1245_));
 sky130_fd_sc_hd__and2_4 _4283_ (.A(_1950_),
    .B(_1954_),
    .X(_1956_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_1947_),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__and4_4 _4285_ (.A(_1943_),
    .B(_1945_),
    .C(_1947_),
    .D(_1956_),
    .X(_1958_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(_1941_),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__and4_1 _4287_ (.A(_1936_),
    .B(_1939_),
    .C(_1941_),
    .D(_1958_),
    .X(_1960_));
 sky130_fd_sc_hd__nand2_1 _4288_ (.A(_1934_),
    .B(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__and4_1 _4289_ (.A(_1929_),
    .B(_1932_),
    .C(_1934_),
    .D(_1960_),
    .X(_1962_));
 sky130_fd_sc_hd__nand2_1 _4290_ (.A(_1927_),
    .B(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__and4_4 _4291_ (.A(_1922_),
    .B(_1925_),
    .C(_1927_),
    .D(_1962_),
    .X(_1964_));
 sky130_fd_sc_hd__and3_1 _4292_ (.A(_1918_),
    .B(_1920_),
    .C(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__and2_4 _4293_ (.A(_1916_),
    .B(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__nand2_4 _4294_ (.A(_1914_),
    .B(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__nor2_2 _4295_ (.A(_1912_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__and2_1 _4296_ (.A(_1908_),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_1906_),
    .B(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__and3_1 _4298_ (.A(_1904_),
    .B(_1906_),
    .C(_1969_),
    .X(_1971_));
 sky130_fd_sc_hd__and2_4 _4299_ (.A(_1901_),
    .B(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__nand2_1 _4300_ (.A(_1899_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__nand2b_1 _4301_ (.A_N(_1973_),
    .B(_1896_),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2b_2 _4302_ (.A_N(_1974_),
    .B(_1893_),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2b_4 _4303_ (.A_N(_1975_),
    .B(_1890_),
    .Y(_1976_));
 sky130_fd_sc_hd__and2b_1 _4304_ (.A_N(_1976_),
    .B(_1887_),
    .X(_1977_));
 sky130_fd_sc_hd__nor2_1 _4305_ (.A(net254),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__nand2_2 _4306_ (.A(_1884_),
    .B(_1977_),
    .Y(_1979_));
 sky130_fd_sc_hd__xnor2_1 _4307_ (.A(_1882_),
    .B(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(net2041),
    .A1(_1980_),
    .S(net247),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _4309_ (.A(_1884_),
    .B(_1977_),
    .X(_1981_));
 sky130_fd_sc_hd__and2_1 _4310_ (.A(net2061),
    .B(net254),
    .X(_1982_));
 sky130_fd_sc_hd__a31o_1 _4311_ (.A1(net245),
    .A2(_1979_),
    .A3(_1981_),
    .B1(_1982_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2b_1 _4312_ (.A_N(_1887_),
    .B(_1976_),
    .Y(_1983_));
 sky130_fd_sc_hd__a22o_1 _4313_ (.A1(net2051),
    .A2(net254),
    .B1(_1978_),
    .B2(_1983_),
    .X(_0320_));
 sky130_fd_sc_hd__and2_1 _4314_ (.A(net2025),
    .B(net254),
    .X(_1984_));
 sky130_fd_sc_hd__nand2b_1 _4315_ (.A_N(_1890_),
    .B(_1975_),
    .Y(_1985_));
 sky130_fd_sc_hd__a31o_1 _4316_ (.A1(net244),
    .A2(_1976_),
    .A3(_1985_),
    .B1(_1984_),
    .X(_0319_));
 sky130_fd_sc_hd__and2_1 _4317_ (.A(net2066),
    .B(net255),
    .X(_1986_));
 sky130_fd_sc_hd__a31o_1 _4318_ (.A1(_1896_),
    .A2(_1899_),
    .A3(_1972_),
    .B1(_1893_),
    .X(_1987_));
 sky130_fd_sc_hd__a31o_1 _4319_ (.A1(net246),
    .A2(_1975_),
    .A3(_1987_),
    .B1(_1986_),
    .X(_0318_));
 sky130_fd_sc_hd__and2_1 _4320_ (.A(net1955),
    .B(net255),
    .X(_1988_));
 sky130_fd_sc_hd__a21o_1 _4321_ (.A1(_1899_),
    .A2(_1972_),
    .B1(_1896_),
    .X(_1989_));
 sky130_fd_sc_hd__a31o_1 _4322_ (.A1(net246),
    .A2(_1974_),
    .A3(_1989_),
    .B1(_1988_),
    .X(_0317_));
 sky130_fd_sc_hd__and2_1 _4323_ (.A(net2036),
    .B(net255),
    .X(_1990_));
 sky130_fd_sc_hd__or2_1 _4324_ (.A(_1899_),
    .B(_1972_),
    .X(_1991_));
 sky130_fd_sc_hd__a31o_1 _4325_ (.A1(net246),
    .A2(_1973_),
    .A3(_1991_),
    .B1(_1990_),
    .X(_0316_));
 sky130_fd_sc_hd__or2_1 _4326_ (.A(_1901_),
    .B(_1971_),
    .X(_1992_));
 sky130_fd_sc_hd__nor2_1 _4327_ (.A(net255),
    .B(_1972_),
    .Y(_1993_));
 sky130_fd_sc_hd__a22o_1 _4328_ (.A1(net2047),
    .A2(net255),
    .B1(_1992_),
    .B2(_1993_),
    .X(_0315_));
 sky130_fd_sc_hd__a31o_1 _4329_ (.A1(_1906_),
    .A2(_1908_),
    .A3(_1968_),
    .B1(_1904_),
    .X(_1994_));
 sky130_fd_sc_hd__nor2_1 _4330_ (.A(net255),
    .B(_1971_),
    .Y(_1995_));
 sky130_fd_sc_hd__a22o_1 _4331_ (.A1(net2073),
    .A2(net255),
    .B1(_1994_),
    .B2(_1995_),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _4332_ (.A(net2060),
    .B(net254),
    .X(_1996_));
 sky130_fd_sc_hd__or2_1 _4333_ (.A(_1906_),
    .B(_1969_),
    .X(_1997_));
 sky130_fd_sc_hd__a31o_1 _4334_ (.A1(net244),
    .A2(_1970_),
    .A3(_1997_),
    .B1(_1996_),
    .X(_0313_));
 sky130_fd_sc_hd__or2_1 _4335_ (.A(_1908_),
    .B(_1968_),
    .X(_1998_));
 sky130_fd_sc_hd__nor2_1 _4336_ (.A(net255),
    .B(_1969_),
    .Y(_1999_));
 sky130_fd_sc_hd__a22o_1 _4337_ (.A1(net2033),
    .A2(net255),
    .B1(_1998_),
    .B2(_1999_),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _4338_ (.A(_1912_),
    .B(_1967_),
    .X(_2000_));
 sky130_fd_sc_hd__nor2_1 _4339_ (.A(_1968_),
    .B(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(net2007),
    .A1(_2001_),
    .S(net246),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _4341_ (.A(net2049),
    .B(net261),
    .X(_2002_));
 sky130_fd_sc_hd__or2_1 _4342_ (.A(_1914_),
    .B(_1966_),
    .X(_2003_));
 sky130_fd_sc_hd__a31o_1 _4343_ (.A1(_1324_),
    .A2(_1967_),
    .A3(_2003_),
    .B1(_2002_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _4344_ (.A(_1916_),
    .B(_1965_),
    .X(_2004_));
 sky130_fd_sc_hd__nor2_1 _4345_ (.A(net259),
    .B(_1966_),
    .Y(_2005_));
 sky130_fd_sc_hd__a22o_1 _4346_ (.A1(net889),
    .A2(net259),
    .B1(_2004_),
    .B2(_2005_),
    .X(_0309_));
 sky130_fd_sc_hd__a21o_1 _4347_ (.A1(_1920_),
    .A2(_1964_),
    .B1(_1918_),
    .X(_2006_));
 sky130_fd_sc_hd__nor2_1 _4348_ (.A(net260),
    .B(_1965_),
    .Y(_2007_));
 sky130_fd_sc_hd__a22o_1 _4349_ (.A1(net2034),
    .A2(net260),
    .B1(_2006_),
    .B2(_2007_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _4350_ (.A(_1920_),
    .B(_1964_),
    .X(_2008_));
 sky130_fd_sc_hd__a21oi_1 _4351_ (.A1(_1920_),
    .A2(_1964_),
    .B1(net259),
    .Y(_2009_));
 sky130_fd_sc_hd__a22o_1 _4352_ (.A1(net2062),
    .A2(net260),
    .B1(_2008_),
    .B2(_2009_),
    .X(_0307_));
 sky130_fd_sc_hd__a31o_1 _4353_ (.A1(_1925_),
    .A2(_1927_),
    .A3(_1962_),
    .B1(_1922_),
    .X(_2010_));
 sky130_fd_sc_hd__nor2_1 _4354_ (.A(net262),
    .B(_1964_),
    .Y(_2011_));
 sky130_fd_sc_hd__a22o_1 _4355_ (.A1(net2083),
    .A2(net262),
    .B1(_2010_),
    .B2(_2011_),
    .X(_0306_));
 sky130_fd_sc_hd__xnor2_1 _4356_ (.A(_1925_),
    .B(_1963_),
    .Y(_2012_));
 sky130_fd_sc_hd__mux2_1 _4357_ (.A0(net2009),
    .A1(_2012_),
    .S(net251),
    .X(_0305_));
 sky130_fd_sc_hd__and2_1 _4358_ (.A(net2027),
    .B(net262),
    .X(_2013_));
 sky130_fd_sc_hd__or2_1 _4359_ (.A(_1927_),
    .B(_1962_),
    .X(_2014_));
 sky130_fd_sc_hd__a31o_1 _4360_ (.A1(net251),
    .A2(_1963_),
    .A3(_2014_),
    .B1(_2013_),
    .X(_0304_));
 sky130_fd_sc_hd__a31o_1 _4361_ (.A1(_1932_),
    .A2(_1934_),
    .A3(_1960_),
    .B1(_1929_),
    .X(_2015_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(net262),
    .B(_1962_),
    .Y(_2016_));
 sky130_fd_sc_hd__a22o_1 _4363_ (.A1(net1741),
    .A2(net262),
    .B1(_2015_),
    .B2(_2016_),
    .X(_0303_));
 sky130_fd_sc_hd__xnor2_1 _4364_ (.A(_1932_),
    .B(_1961_),
    .Y(_2017_));
 sky130_fd_sc_hd__mux2_1 _4365_ (.A0(net2065),
    .A1(_2017_),
    .S(net249),
    .X(_0302_));
 sky130_fd_sc_hd__and2_1 _4366_ (.A(net2043),
    .B(net259),
    .X(_2018_));
 sky130_fd_sc_hd__or2_1 _4367_ (.A(_1934_),
    .B(_1960_),
    .X(_2019_));
 sky130_fd_sc_hd__a31o_1 _4368_ (.A1(net251),
    .A2(_1961_),
    .A3(_2019_),
    .B1(_2018_),
    .X(_0301_));
 sky130_fd_sc_hd__a31o_1 _4369_ (.A1(_1939_),
    .A2(_1941_),
    .A3(_1958_),
    .B1(_1936_),
    .X(_2020_));
 sky130_fd_sc_hd__nor2_1 _4370_ (.A(net262),
    .B(_1960_),
    .Y(_2021_));
 sky130_fd_sc_hd__a22o_1 _4371_ (.A1(net2016),
    .A2(net262),
    .B1(_2020_),
    .B2(_2021_),
    .X(_0300_));
 sky130_fd_sc_hd__xnor2_1 _4372_ (.A(_1939_),
    .B(_1959_),
    .Y(_2022_));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(net2017),
    .A1(_2022_),
    .S(net249),
    .X(_0299_));
 sky130_fd_sc_hd__and2_1 _4374_ (.A(net949),
    .B(net259),
    .X(_2023_));
 sky130_fd_sc_hd__or2_1 _4375_ (.A(_1941_),
    .B(_1958_),
    .X(_2024_));
 sky130_fd_sc_hd__a31o_1 _4376_ (.A1(net249),
    .A2(_1959_),
    .A3(_2024_),
    .B1(_2023_),
    .X(_0298_));
 sky130_fd_sc_hd__a31o_1 _4377_ (.A1(_1945_),
    .A2(_1947_),
    .A3(_1956_),
    .B1(_1943_),
    .X(_2025_));
 sky130_fd_sc_hd__or3b_1 _4378_ (.A(net262),
    .B(_1958_),
    .C_N(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__a21bo_1 _4379_ (.A1(net1998),
    .A2(net262),
    .B1_N(_2026_),
    .X(_0297_));
 sky130_fd_sc_hd__xnor2_1 _4380_ (.A(_1945_),
    .B(_1957_),
    .Y(_2027_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(net2008),
    .A1(_2027_),
    .S(net251),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_1 _4382_ (.A(_1947_),
    .B(_1956_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _4383_ (.A(net251),
    .B(_1957_),
    .Y(_2029_));
 sky130_fd_sc_hd__a2bb2o_1 _4384_ (.A1_N(_2028_),
    .A2_N(_2029_),
    .B1(net2015),
    .B2(net262),
    .X(_0295_));
 sky130_fd_sc_hd__nor2_1 _4385_ (.A(_1950_),
    .B(_1954_),
    .Y(_2030_));
 sky130_fd_sc_hd__or2_1 _4386_ (.A(net263),
    .B(_1956_),
    .X(_2031_));
 sky130_fd_sc_hd__a2bb2o_1 _4387_ (.A1_N(_2030_),
    .A2_N(_2031_),
    .B1(net2040),
    .B2(net263),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _4388_ (.A1(net2082),
    .A2(net264),
    .B1(_1955_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_2 _4389_ (.A(net2037),
    .B(net2076),
    .Y(_2032_));
 sky130_fd_sc_hd__or4_4 _4390_ (.A(net2170),
    .B(net919),
    .C(net2037),
    .D(net2076),
    .X(_2033_));
 sky130_fd_sc_hd__and4b_2 _4391_ (.A_N(net919),
    .B(net2076),
    .C(net2170),
    .D(net2029),
    .X(_2034_));
 sky130_fd_sc_hd__or4b_4 _4392_ (.A(_1280_),
    .B(_1281_),
    .C(net919),
    .D_N(net2076),
    .X(_2035_));
 sky130_fd_sc_hd__and4_4 _4393_ (.A(_1280_),
    .B(net919),
    .C(_1282_),
    .D(net2076),
    .X(_2036_));
 sky130_fd_sc_hd__or4bb_4 _4394_ (.A(net2237),
    .B(net2037),
    .C_N(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .D_N(net919),
    .X(_2037_));
 sky130_fd_sc_hd__or2_1 _4395_ (.A(_2034_),
    .B(_2036_),
    .X(_2038_));
 sky130_fd_sc_hd__o211a_1 _4396_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .A2(_2037_),
    .B1(_2035_),
    .C1(_2033_),
    .X(_3562_));
 sky130_fd_sc_hd__mux4_1 _4397_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net424),
    .S1(net414),
    .X(_2039_));
 sky130_fd_sc_hd__mux4_1 _4398_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net424),
    .S1(net414),
    .X(_2040_));
 sky130_fd_sc_hd__mux2_1 _4399_ (.A0(_2039_),
    .A1(_2040_),
    .S(net403),
    .X(_2041_));
 sky130_fd_sc_hd__mux4_1 _4400_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net422),
    .S1(net411),
    .X(_2042_));
 sky130_fd_sc_hd__mux4_1 _4401_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net422),
    .S1(net411),
    .X(_2043_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(_2043_),
    .A1(_2042_),
    .S(net403),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _4403_ (.A0(_2044_),
    .A1(_2041_),
    .S(net398),
    .X(_0032_));
 sky130_fd_sc_hd__mux4_1 _4404_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net424),
    .S1(net414),
    .X(_2045_));
 sky130_fd_sc_hd__mux4_1 _4405_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net422),
    .S1(net411),
    .X(_2046_));
 sky130_fd_sc_hd__mux2_1 _4406_ (.A0(_2045_),
    .A1(_2046_),
    .S(net403),
    .X(_2047_));
 sky130_fd_sc_hd__mux4_1 _4407_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net422),
    .S1(net410),
    .X(_2048_));
 sky130_fd_sc_hd__mux4_1 _4408_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net421),
    .S1(net410),
    .X(_2049_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(_2049_),
    .A1(_2048_),
    .S(net402),
    .X(_2050_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(_2050_),
    .A1(_2047_),
    .S(net398),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_1 _4411_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net421),
    .S1(net410),
    .X(_2051_));
 sky130_fd_sc_hd__mux4_1 _4412_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net424),
    .S1(net414),
    .X(_2052_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(_2051_),
    .A1(_2052_),
    .S(net403),
    .X(_2053_));
 sky130_fd_sc_hd__mux4_1 _4414_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net421),
    .S1(net411),
    .X(_2054_));
 sky130_fd_sc_hd__mux4_1 _4415_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net421),
    .S1(net411),
    .X(_2055_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(_2055_),
    .A1(_2054_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(_2056_));
 sky130_fd_sc_hd__mux2_1 _4417_ (.A0(_2056_),
    .A1(_2053_),
    .S(net398),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_1 _4418_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net424),
    .S1(net414),
    .X(_2057_));
 sky130_fd_sc_hd__mux4_1 _4419_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net424),
    .S1(net414),
    .X(_2058_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(_2057_),
    .A1(_2058_),
    .S(net404),
    .X(_2059_));
 sky130_fd_sc_hd__mux4_1 _4421_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net424),
    .S1(net413),
    .X(_2060_));
 sky130_fd_sc_hd__mux4_1 _4422_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net424),
    .S1(net413),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(_2061_),
    .A1(_2060_),
    .S(net404),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_1 _4424_ (.A0(_2062_),
    .A1(_2059_),
    .S(net398),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_1 _4425_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net423),
    .S1(net412),
    .X(_2063_));
 sky130_fd_sc_hd__mux4_1 _4426_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net423),
    .S1(net412),
    .X(_2064_));
 sky130_fd_sc_hd__mux2_1 _4427_ (.A0(_2063_),
    .A1(_2064_),
    .S(net403),
    .X(_2065_));
 sky130_fd_sc_hd__mux4_1 _4428_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net423),
    .S1(net412),
    .X(_2066_));
 sky130_fd_sc_hd__mux4_1 _4429_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net423),
    .S1(net412),
    .X(_2067_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(_2067_),
    .A1(_2066_),
    .S(net403),
    .X(_2068_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(_2068_),
    .A1(_2065_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _4432_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net423),
    .S1(net412),
    .X(_2069_));
 sky130_fd_sc_hd__mux4_1 _4433_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net423),
    .S1(net414),
    .X(_2070_));
 sky130_fd_sc_hd__mux2_1 _4434_ (.A0(_2069_),
    .A1(_2070_),
    .S(net403),
    .X(_2071_));
 sky130_fd_sc_hd__mux4_1 _4435_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net425),
    .S1(net412),
    .X(_2072_));
 sky130_fd_sc_hd__mux4_1 _4436_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net425),
    .S1(net412),
    .X(_2073_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(_2073_),
    .A1(_2072_),
    .S(net404),
    .X(_2074_));
 sky130_fd_sc_hd__mux2_1 _4438_ (.A0(_2074_),
    .A1(_2071_),
    .S(net398),
    .X(_0059_));
 sky130_fd_sc_hd__mux4_1 _4439_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net419),
    .S1(net408),
    .X(_2075_));
 sky130_fd_sc_hd__mux4_1 _4440_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net420),
    .S1(net409),
    .X(_2076_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(_2075_),
    .A1(_2076_),
    .S(net401),
    .X(_2077_));
 sky130_fd_sc_hd__mux4_1 _4442_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net420),
    .S1(net409),
    .X(_2078_));
 sky130_fd_sc_hd__mux4_1 _4443_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net419),
    .S1(net408),
    .X(_2079_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(_2079_),
    .A1(_2078_),
    .S(net401),
    .X(_2080_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(_2080_),
    .A1(_2077_),
    .S(net399),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _4446_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net421),
    .S1(net410),
    .X(_2081_));
 sky130_fd_sc_hd__mux4_1 _4447_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net421),
    .S1(net410),
    .X(_2082_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(_2081_),
    .A1(_2082_),
    .S(net402),
    .X(_2083_));
 sky130_fd_sc_hd__mux4_1 _4449_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net421),
    .S1(net410),
    .X(_2084_));
 sky130_fd_sc_hd__mux4_1 _4450_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net421),
    .S1(net410),
    .X(_2085_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(_2085_),
    .A1(_2084_),
    .S(net402),
    .X(_2086_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(_2086_),
    .A1(_2083_),
    .S(net398),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_1 _4453_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net422),
    .S1(net410),
    .X(_2087_));
 sky130_fd_sc_hd__mux4_1 _4454_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net422),
    .S1(net410),
    .X(_2088_));
 sky130_fd_sc_hd__mux2_1 _4455_ (.A0(_2087_),
    .A1(_2088_),
    .S(net402),
    .X(_2089_));
 sky130_fd_sc_hd__mux4_1 _4456_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(net420),
    .S1(net408),
    .X(_2090_));
 sky130_fd_sc_hd__mux4_1 _4457_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net420),
    .S1(net409),
    .X(_2091_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(_2091_),
    .A1(_2090_),
    .S(net402),
    .X(_2092_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(_2092_),
    .A1(_2089_),
    .S(net398),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_1 _4460_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net424),
    .S1(net413),
    .X(_2093_));
 sky130_fd_sc_hd__mux4_1 _4461_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net424),
    .S1(net413),
    .X(_2094_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(_2093_),
    .A1(_2094_),
    .S(net404),
    .X(_2095_));
 sky130_fd_sc_hd__mux4_1 _4463_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net424),
    .S1(net413),
    .X(_2096_));
 sky130_fd_sc_hd__mux4_1 _4464_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net424),
    .S1(net413),
    .X(_2097_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(_2097_),
    .A1(_2096_),
    .S(net404),
    .X(_2098_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(_2098_),
    .A1(_2095_),
    .S(net398),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _4467_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(net419),
    .S1(net408),
    .X(_2099_));
 sky130_fd_sc_hd__mux4_1 _4468_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(net419),
    .S1(net409),
    .X(_2100_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(_2099_),
    .A1(_2100_),
    .S(net402),
    .X(_2101_));
 sky130_fd_sc_hd__mux4_1 _4470_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net419),
    .S1(net408),
    .X(_2102_));
 sky130_fd_sc_hd__mux4_1 _4471_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net419),
    .S1(net408),
    .X(_2103_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(_2103_),
    .A1(_2102_),
    .S(net402),
    .X(_2104_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(_2104_),
    .A1(_2101_),
    .S(net398),
    .X(_0033_));
 sky130_fd_sc_hd__mux4_1 _4474_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net418),
    .S1(net405),
    .X(_2105_));
 sky130_fd_sc_hd__mux4_1 _4475_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net418),
    .S1(net407),
    .X(_2106_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(_2105_),
    .A1(_2106_),
    .S(net400),
    .X(_2107_));
 sky130_fd_sc_hd__mux4_1 _4477_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net418),
    .S1(net405),
    .X(_2108_));
 sky130_fd_sc_hd__mux4_1 _4478_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net418),
    .S1(net405),
    .X(_2109_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(_2109_),
    .A1(_2108_),
    .S(net400),
    .X(_2110_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(_2110_),
    .A1(_2107_),
    .S(net399),
    .X(_0034_));
 sky130_fd_sc_hd__mux4_1 _4481_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net425),
    .S1(net412),
    .X(_2111_));
 sky130_fd_sc_hd__mux4_1 _4482_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net425),
    .S1(net412),
    .X(_2112_));
 sky130_fd_sc_hd__mux2_1 _4483_ (.A0(_2111_),
    .A1(_2112_),
    .S(net403),
    .X(_2113_));
 sky130_fd_sc_hd__mux4_1 _4484_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net425),
    .S1(net412),
    .X(_2114_));
 sky130_fd_sc_hd__mux4_1 _4485_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net425),
    .S1(net412),
    .X(_2115_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(_2115_),
    .A1(_2114_),
    .S(net403),
    .X(_2116_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(_2116_),
    .A1(_2113_),
    .S(net398),
    .X(_0035_));
 sky130_fd_sc_hd__mux4_1 _4488_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net419),
    .S1(net408),
    .X(_2117_));
 sky130_fd_sc_hd__mux4_1 _4489_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net419),
    .S1(net408),
    .X(_2118_));
 sky130_fd_sc_hd__mux2_1 _4490_ (.A0(_2117_),
    .A1(_2118_),
    .S(net401),
    .X(_2119_));
 sky130_fd_sc_hd__mux4_1 _4491_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net419),
    .S1(net408),
    .X(_2120_));
 sky130_fd_sc_hd__mux4_1 _4492_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net419),
    .S1(net408),
    .X(_2121_));
 sky130_fd_sc_hd__mux2_1 _4493_ (.A0(_2121_),
    .A1(_2120_),
    .S(net401),
    .X(_2122_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(_2122_),
    .A1(_2119_),
    .S(net399),
    .X(_0036_));
 sky130_fd_sc_hd__mux4_1 _4495_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net423),
    .S1(net414),
    .X(_2123_));
 sky130_fd_sc_hd__mux4_1 _4496_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net423),
    .S1(net414),
    .X(_2124_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(_2123_),
    .A1(_2124_),
    .S(net403),
    .X(_2125_));
 sky130_fd_sc_hd__mux4_1 _4498_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net423),
    .S1(net414),
    .X(_2126_));
 sky130_fd_sc_hd__mux4_1 _4499_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net423),
    .S1(net414),
    .X(_2127_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(_2127_),
    .A1(_2126_),
    .S(net403),
    .X(_2128_));
 sky130_fd_sc_hd__mux2_1 _4501_ (.A0(_2128_),
    .A1(_2125_),
    .S(net398),
    .X(_0037_));
 sky130_fd_sc_hd__mux4_1 _4502_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net422),
    .S1(net411),
    .X(_2129_));
 sky130_fd_sc_hd__mux4_1 _4503_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net422),
    .S1(net411),
    .X(_2130_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(_2129_),
    .A1(_2130_),
    .S(net403),
    .X(_2131_));
 sky130_fd_sc_hd__mux4_1 _4505_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net423),
    .S1(net414),
    .X(_2132_));
 sky130_fd_sc_hd__mux4_1 _4506_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net422),
    .S1(net411),
    .X(_2133_));
 sky130_fd_sc_hd__mux2_1 _4507_ (.A0(_2133_),
    .A1(_2132_),
    .S(net403),
    .X(_2134_));
 sky130_fd_sc_hd__mux2_1 _4508_ (.A0(_2134_),
    .A1(_2131_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _4509_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net420),
    .S1(net409),
    .X(_2135_));
 sky130_fd_sc_hd__mux4_1 _4510_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net421),
    .S1(net410),
    .X(_2136_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(_2135_),
    .A1(_2136_),
    .S(net402),
    .X(_2137_));
 sky130_fd_sc_hd__mux4_1 _4512_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net419),
    .S1(net409),
    .X(_2138_));
 sky130_fd_sc_hd__mux4_1 _4513_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net421),
    .S1(net410),
    .X(_2139_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(_2139_),
    .A1(_2138_),
    .S(net402),
    .X(_2140_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(_2140_),
    .A1(_2137_),
    .S(net398),
    .X(_0039_));
 sky130_fd_sc_hd__mux4_1 _4516_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net421),
    .S1(net411),
    .X(_2141_));
 sky130_fd_sc_hd__mux4_1 _4517_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net421),
    .S1(net411),
    .X(_2142_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(_2141_),
    .A1(_2142_),
    .S(net402),
    .X(_2143_));
 sky130_fd_sc_hd__mux4_1 _4519_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net422),
    .S1(net411),
    .X(_2144_));
 sky130_fd_sc_hd__mux4_1 _4520_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net422),
    .S1(net411),
    .X(_2145_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(_2145_),
    .A1(_2144_),
    .S(net402),
    .X(_2146_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(_2146_),
    .A1(_2143_),
    .S(net398),
    .X(_0040_));
 sky130_fd_sc_hd__mux4_1 _4523_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net424),
    .S1(net412),
    .X(_2147_));
 sky130_fd_sc_hd__mux4_1 _4524_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net423),
    .S1(net412),
    .X(_2148_));
 sky130_fd_sc_hd__mux2_1 _4525_ (.A0(_2147_),
    .A1(_2148_),
    .S(net404),
    .X(_2149_));
 sky130_fd_sc_hd__mux4_1 _4526_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net423),
    .S1(net412),
    .X(_2150_));
 sky130_fd_sc_hd__mux4_1 _4527_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net423),
    .S1(net412),
    .X(_2151_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(_2151_),
    .A1(_2150_),
    .S(net404),
    .X(_2152_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(_2152_),
    .A1(_2149_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0041_));
 sky130_fd_sc_hd__mux4_1 _4530_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net419),
    .S1(net408),
    .X(_2153_));
 sky130_fd_sc_hd__mux4_1 _4531_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net419),
    .S1(net408),
    .X(_2154_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(_2153_),
    .A1(_2154_),
    .S(net400),
    .X(_2155_));
 sky130_fd_sc_hd__mux4_1 _4533_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net419),
    .S1(net408),
    .X(_2156_));
 sky130_fd_sc_hd__mux4_1 _4534_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net419),
    .S1(net408),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(_2157_),
    .A1(_2156_),
    .S(net400),
    .X(_2158_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(_2158_),
    .A1(_2155_),
    .S(net399),
    .X(_0042_));
 sky130_fd_sc_hd__mux4_1 _4537_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net418),
    .S1(net407),
    .X(_2159_));
 sky130_fd_sc_hd__mux4_1 _4538_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net418),
    .S1(net407),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(_2159_),
    .A1(_2160_),
    .S(net401),
    .X(_2161_));
 sky130_fd_sc_hd__mux4_1 _4540_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net417),
    .S1(net407),
    .X(_2162_));
 sky130_fd_sc_hd__mux4_1 _4541_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net418),
    .S1(net407),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(_2163_),
    .A1(_2162_),
    .S(net401),
    .X(_2164_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(_2164_),
    .A1(_2161_),
    .S(net399),
    .X(_0044_));
 sky130_fd_sc_hd__mux4_1 _4544_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net417),
    .S1(net407),
    .X(_2165_));
 sky130_fd_sc_hd__mux4_1 _4545_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net417),
    .S1(net407),
    .X(_2166_));
 sky130_fd_sc_hd__mux2_1 _4546_ (.A0(_2165_),
    .A1(_2166_),
    .S(net401),
    .X(_2167_));
 sky130_fd_sc_hd__mux4_1 _4547_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net417),
    .S1(net407),
    .X(_2168_));
 sky130_fd_sc_hd__mux4_1 _4548_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net417),
    .S1(net407),
    .X(_2169_));
 sky130_fd_sc_hd__mux2_1 _4549_ (.A0(_2169_),
    .A1(_2168_),
    .S(net401),
    .X(_2170_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(_2170_),
    .A1(_2167_),
    .S(net399),
    .X(_0045_));
 sky130_fd_sc_hd__mux4_1 _4551_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net421),
    .S1(net410),
    .X(_2171_));
 sky130_fd_sc_hd__mux4_1 _4552_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net421),
    .S1(net410),
    .X(_2172_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(_2171_),
    .A1(_2172_),
    .S(net402),
    .X(_2173_));
 sky130_fd_sc_hd__mux4_1 _4554_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net421),
    .S1(net410),
    .X(_2174_));
 sky130_fd_sc_hd__mux4_1 _4555_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net421),
    .S1(net410),
    .X(_2175_));
 sky130_fd_sc_hd__mux2_1 _4556_ (.A0(_2175_),
    .A1(_2174_),
    .S(net402),
    .X(_2176_));
 sky130_fd_sc_hd__mux2_1 _4557_ (.A0(_2176_),
    .A1(_2173_),
    .S(net398),
    .X(_0046_));
 sky130_fd_sc_hd__mux4_1 _4558_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net416),
    .S1(net405),
    .X(_2177_));
 sky130_fd_sc_hd__mux4_1 _4559_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net416),
    .S1(net405),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_1 _4560_ (.A0(_2177_),
    .A1(_2178_),
    .S(net400),
    .X(_2179_));
 sky130_fd_sc_hd__mux4_1 _4561_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net416),
    .S1(net406),
    .X(_2180_));
 sky130_fd_sc_hd__mux4_1 _4562_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net416),
    .S1(net406),
    .X(_2181_));
 sky130_fd_sc_hd__mux2_1 _4563_ (.A0(_2181_),
    .A1(_2180_),
    .S(net400),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _4564_ (.A0(_2182_),
    .A1(_2179_),
    .S(net399),
    .X(_0047_));
 sky130_fd_sc_hd__mux4_1 _4565_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net425),
    .S1(net413),
    .X(_2183_));
 sky130_fd_sc_hd__mux4_1 _4566_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net424),
    .S1(net412),
    .X(_2184_));
 sky130_fd_sc_hd__mux2_1 _4567_ (.A0(_2183_),
    .A1(_2184_),
    .S(net404),
    .X(_2185_));
 sky130_fd_sc_hd__mux4_1 _4568_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net425),
    .S1(net413),
    .X(_2186_));
 sky130_fd_sc_hd__mux4_1 _4569_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net424),
    .S1(net413),
    .X(_2187_));
 sky130_fd_sc_hd__mux2_1 _4570_ (.A0(_2187_),
    .A1(_2186_),
    .S(net404),
    .X(_2188_));
 sky130_fd_sc_hd__mux2_1 _4571_ (.A0(_2188_),
    .A1(_2185_),
    .S(net398),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _4572_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net416),
    .S1(net405),
    .X(_2189_));
 sky130_fd_sc_hd__mux4_1 _4573_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net416),
    .S1(net405),
    .X(_2190_));
 sky130_fd_sc_hd__mux2_1 _4574_ (.A0(_2189_),
    .A1(_2190_),
    .S(net400),
    .X(_2191_));
 sky130_fd_sc_hd__mux4_1 _4575_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net416),
    .S1(net406),
    .X(_2192_));
 sky130_fd_sc_hd__mux4_1 _4576_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net416),
    .S1(net406),
    .X(_2193_));
 sky130_fd_sc_hd__mux2_1 _4577_ (.A0(_2193_),
    .A1(_2192_),
    .S(net400),
    .X(_2194_));
 sky130_fd_sc_hd__mux2_1 _4578_ (.A0(_2194_),
    .A1(_2191_),
    .S(net399),
    .X(_0049_));
 sky130_fd_sc_hd__mux4_1 _4579_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2195_));
 sky130_fd_sc_hd__mux4_1 _4580_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2196_));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(_2195_),
    .A1(_2196_),
    .S(net400),
    .X(_2197_));
 sky130_fd_sc_hd__mux4_1 _4582_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2198_));
 sky130_fd_sc_hd__mux4_1 _4583_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2199_));
 sky130_fd_sc_hd__mux2_1 _4584_ (.A0(_2199_),
    .A1(_2198_),
    .S(net400),
    .X(_2200_));
 sky130_fd_sc_hd__mux2_1 _4585_ (.A0(_2200_),
    .A1(_2197_),
    .S(net399),
    .X(_0050_));
 sky130_fd_sc_hd__mux4_1 _4586_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net420),
    .S1(net409),
    .X(_2201_));
 sky130_fd_sc_hd__mux4_1 _4587_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net420),
    .S1(net409),
    .X(_2202_));
 sky130_fd_sc_hd__mux2_1 _4588_ (.A0(_2201_),
    .A1(_2202_),
    .S(net402),
    .X(_2203_));
 sky130_fd_sc_hd__mux4_1 _4589_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net420),
    .S1(net409),
    .X(_2204_));
 sky130_fd_sc_hd__mux4_1 _4590_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net420),
    .S1(net409),
    .X(_2205_));
 sky130_fd_sc_hd__mux2_1 _4591_ (.A0(_2205_),
    .A1(_2204_),
    .S(net402),
    .X(_2206_));
 sky130_fd_sc_hd__mux2_1 _4592_ (.A0(_2206_),
    .A1(_2203_),
    .S(net399),
    .X(_0051_));
 sky130_fd_sc_hd__mux4_1 _4593_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net418),
    .S1(net405),
    .X(_2207_));
 sky130_fd_sc_hd__mux4_1 _4594_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net418),
    .S1(net405),
    .X(_2208_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(_2207_),
    .A1(_2208_),
    .S(net400),
    .X(_2209_));
 sky130_fd_sc_hd__mux4_1 _4596_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net418),
    .S1(net405),
    .X(_2210_));
 sky130_fd_sc_hd__mux4_1 _4597_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net418),
    .S1(net405),
    .X(_2211_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(_2211_),
    .A1(_2210_),
    .S(net400),
    .X(_2212_));
 sky130_fd_sc_hd__mux2_1 _4599_ (.A0(_2212_),
    .A1(_2209_),
    .S(net399),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _4600_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net418),
    .S1(net405),
    .X(_2213_));
 sky130_fd_sc_hd__mux4_1 _4601_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net418),
    .S1(net405),
    .X(_2214_));
 sky130_fd_sc_hd__mux2_1 _4602_ (.A0(_2213_),
    .A1(_2214_),
    .S(net400),
    .X(_2215_));
 sky130_fd_sc_hd__mux4_1 _4603_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net418),
    .S1(net405),
    .X(_2216_));
 sky130_fd_sc_hd__mux4_1 _4604_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net418),
    .S1(net405),
    .X(_2217_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(_2217_),
    .A1(_2216_),
    .S(net400),
    .X(_2218_));
 sky130_fd_sc_hd__mux2_1 _4606_ (.A0(_2218_),
    .A1(_2215_),
    .S(net399),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_1 _4607_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net417),
    .S1(net407),
    .X(_2219_));
 sky130_fd_sc_hd__mux4_1 _4608_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net417),
    .S1(net407),
    .X(_2220_));
 sky130_fd_sc_hd__mux2_1 _4609_ (.A0(_2219_),
    .A1(_2220_),
    .S(net401),
    .X(_2221_));
 sky130_fd_sc_hd__mux4_1 _4610_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net417),
    .S1(net407),
    .X(_2222_));
 sky130_fd_sc_hd__mux4_1 _4611_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net419),
    .S1(net408),
    .X(_2223_));
 sky130_fd_sc_hd__mux2_1 _4612_ (.A0(_2223_),
    .A1(_2222_),
    .S(net401),
    .X(_2224_));
 sky130_fd_sc_hd__mux2_1 _4613_ (.A0(_2224_),
    .A1(_2221_),
    .S(net399),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _4614_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net416),
    .S1(net407),
    .X(_2225_));
 sky130_fd_sc_hd__mux4_1 _4615_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net416),
    .S1(net407),
    .X(_2226_));
 sky130_fd_sc_hd__mux2_1 _4616_ (.A0(_2225_),
    .A1(_2226_),
    .S(net400),
    .X(_2227_));
 sky130_fd_sc_hd__mux4_1 _4617_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net416),
    .S1(net415),
    .X(_2228_));
 sky130_fd_sc_hd__mux4_1 _4618_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net416),
    .S1(net405),
    .X(_2229_));
 sky130_fd_sc_hd__mux2_1 _4619_ (.A0(_2229_),
    .A1(_2228_),
    .S(net401),
    .X(_2230_));
 sky130_fd_sc_hd__mux2_1 _4620_ (.A0(_2230_),
    .A1(_2227_),
    .S(net399),
    .X(_0056_));
 sky130_fd_sc_hd__mux4_1 _4621_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net395),
    .S1(net385),
    .X(_2231_));
 sky130_fd_sc_hd__mux4_1 _4622_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net395),
    .S1(net385),
    .X(_2232_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(_2231_),
    .A1(_2232_),
    .S(net374),
    .X(_2233_));
 sky130_fd_sc_hd__mux4_1 _4624_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net393),
    .S1(net382),
    .X(_2234_));
 sky130_fd_sc_hd__mux4_1 _4625_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net393),
    .S1(net382),
    .X(_2235_));
 sky130_fd_sc_hd__mux2_1 _4626_ (.A0(_2235_),
    .A1(_2234_),
    .S(net373),
    .X(_2236_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(_2236_),
    .A1(_2233_),
    .S(net370),
    .X(_0000_));
 sky130_fd_sc_hd__mux4_1 _4628_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net395),
    .S1(net385),
    .X(_2237_));
 sky130_fd_sc_hd__mux4_1 _4629_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net393),
    .S1(net382),
    .X(_2238_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(_2237_),
    .A1(_2238_),
    .S(net375),
    .X(_2239_));
 sky130_fd_sc_hd__mux4_1 _4631_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net393),
    .S1(net381),
    .X(_2240_));
 sky130_fd_sc_hd__mux4_1 _4632_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net392),
    .S1(net381),
    .X(_2241_));
 sky130_fd_sc_hd__mux2_1 _4633_ (.A0(_2241_),
    .A1(_2240_),
    .S(net373),
    .X(_2242_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(_2242_),
    .A1(_2239_),
    .S(net369),
    .X(_0011_));
 sky130_fd_sc_hd__mux4_1 _4635_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net393),
    .S1(net382),
    .X(_2243_));
 sky130_fd_sc_hd__mux4_1 _4636_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net395),
    .S1(net385),
    .X(_2244_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(_2243_),
    .A1(_2244_),
    .S(net373),
    .X(_2245_));
 sky130_fd_sc_hd__mux4_1 _4638_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net392),
    .S1(net382),
    .X(_2246_));
 sky130_fd_sc_hd__mux4_1 _4639_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net393),
    .S1(net381),
    .X(_2247_));
 sky130_fd_sc_hd__mux2_1 _4640_ (.A0(_2247_),
    .A1(_2246_),
    .S(net373),
    .X(_2248_));
 sky130_fd_sc_hd__mux2_1 _4641_ (.A0(_2248_),
    .A1(_2245_),
    .S(net369),
    .X(_0022_));
 sky130_fd_sc_hd__mux4_1 _4642_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net395),
    .S1(net385),
    .X(_2249_));
 sky130_fd_sc_hd__mux4_1 _4643_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net395),
    .S1(net385),
    .X(_2250_));
 sky130_fd_sc_hd__mux2_1 _4644_ (.A0(_2249_),
    .A1(_2250_),
    .S(net374),
    .X(_2251_));
 sky130_fd_sc_hd__mux4_1 _4645_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net394),
    .S1(net384),
    .X(_2252_));
 sky130_fd_sc_hd__mux4_1 _4646_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net394),
    .S1(net384),
    .X(_2253_));
 sky130_fd_sc_hd__mux2_1 _4647_ (.A0(_2253_),
    .A1(_2252_),
    .S(net375),
    .X(_2254_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(_2254_),
    .A1(_2251_),
    .S(net370),
    .X(_0025_));
 sky130_fd_sc_hd__mux4_1 _4649_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net394),
    .S1(net383),
    .X(_2255_));
 sky130_fd_sc_hd__mux4_1 _4650_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net394),
    .S1(net383),
    .X(_2256_));
 sky130_fd_sc_hd__mux2_1 _4651_ (.A0(_2255_),
    .A1(_2256_),
    .S(net374),
    .X(_2257_));
 sky130_fd_sc_hd__mux4_1 _4652_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net396),
    .S1(net383),
    .X(_2258_));
 sky130_fd_sc_hd__mux4_1 _4653_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net396),
    .S1(net383),
    .X(_2259_));
 sky130_fd_sc_hd__mux2_1 _4654_ (.A0(_2259_),
    .A1(_2258_),
    .S(net375),
    .X(_2260_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(_2260_),
    .A1(_2257_),
    .S(net369),
    .X(_0026_));
 sky130_fd_sc_hd__mux4_1 _4656_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net396),
    .S1(net383),
    .X(_2261_));
 sky130_fd_sc_hd__mux4_1 _4657_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net396),
    .S1(net385),
    .X(_2262_));
 sky130_fd_sc_hd__mux2_1 _4658_ (.A0(_2261_),
    .A1(_2262_),
    .S(net375),
    .X(_2263_));
 sky130_fd_sc_hd__mux4_1 _4659_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net396),
    .S1(net383),
    .X(_2264_));
 sky130_fd_sc_hd__mux4_1 _4660_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net396),
    .S1(net383),
    .X(_2265_));
 sky130_fd_sc_hd__mux2_1 _4661_ (.A0(_2265_),
    .A1(_2264_),
    .S(net374),
    .X(_2266_));
 sky130_fd_sc_hd__mux2_1 _4662_ (.A0(_2266_),
    .A1(_2263_),
    .S(net369),
    .X(_0027_));
 sky130_fd_sc_hd__mux4_1 _4663_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net390),
    .S1(net379),
    .X(_2267_));
 sky130_fd_sc_hd__mux4_1 _4664_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net391),
    .S1(net380),
    .X(_2268_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(_2267_),
    .A1(_2268_),
    .S(net372),
    .X(_2269_));
 sky130_fd_sc_hd__mux4_1 _4666_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net390),
    .S1(net380),
    .X(_2270_));
 sky130_fd_sc_hd__mux4_1 _4667_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net390),
    .S1(net379),
    .X(_2271_));
 sky130_fd_sc_hd__mux2_1 _4668_ (.A0(_2271_),
    .A1(_2270_),
    .S(net372),
    .X(_2272_));
 sky130_fd_sc_hd__mux2_1 _4669_ (.A0(_2272_),
    .A1(_2269_),
    .S(net368),
    .X(_0028_));
 sky130_fd_sc_hd__mux4_1 _4670_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net392),
    .S1(net381),
    .X(_2273_));
 sky130_fd_sc_hd__mux4_1 _4671_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net392),
    .S1(net381),
    .X(_2274_));
 sky130_fd_sc_hd__mux2_1 _4672_ (.A0(_2273_),
    .A1(_2274_),
    .S(net373),
    .X(_2275_));
 sky130_fd_sc_hd__mux4_1 _4673_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net392),
    .S1(net381),
    .X(_2276_));
 sky130_fd_sc_hd__mux4_1 _4674_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net392),
    .S1(net381),
    .X(_2277_));
 sky130_fd_sc_hd__mux2_1 _4675_ (.A0(_2277_),
    .A1(_2276_),
    .S(net373),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(_2278_),
    .A1(_2275_),
    .S(net369),
    .X(_0029_));
 sky130_fd_sc_hd__mux4_1 _4677_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net392),
    .S1(net381),
    .X(_2279_));
 sky130_fd_sc_hd__mux4_1 _4678_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net392),
    .S1(net381),
    .X(_2280_));
 sky130_fd_sc_hd__mux2_1 _4679_ (.A0(_2279_),
    .A1(_2280_),
    .S(net373),
    .X(_2281_));
 sky130_fd_sc_hd__mux4_1 _4680_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(net390),
    .S1(net379),
    .X(_2282_));
 sky130_fd_sc_hd__mux4_1 _4681_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net390),
    .S1(net380),
    .X(_2283_));
 sky130_fd_sc_hd__mux2_1 _4682_ (.A0(_2283_),
    .A1(_2282_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(_2284_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(_2284_),
    .A1(_2281_),
    .S(net370),
    .X(_0030_));
 sky130_fd_sc_hd__mux4_1 _4684_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net394),
    .S1(net384),
    .X(_2285_));
 sky130_fd_sc_hd__mux4_1 _4685_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net394),
    .S1(net384),
    .X(_2286_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(_2285_),
    .A1(_2286_),
    .S(net375),
    .X(_2287_));
 sky130_fd_sc_hd__mux4_1 _4687_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net394),
    .S1(net384),
    .X(_2288_));
 sky130_fd_sc_hd__mux4_1 _4688_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net394),
    .S1(net384),
    .X(_2289_));
 sky130_fd_sc_hd__mux2_1 _4689_ (.A0(_2289_),
    .A1(_2288_),
    .S(net375),
    .X(_2290_));
 sky130_fd_sc_hd__mux2_1 _4690_ (.A0(_2290_),
    .A1(_2287_),
    .S(net369),
    .X(_0031_));
 sky130_fd_sc_hd__mux4_1 _4691_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(net391),
    .S1(net379),
    .X(_2291_));
 sky130_fd_sc_hd__mux4_1 _4692_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(net391),
    .S1(net380),
    .X(_2292_));
 sky130_fd_sc_hd__mux2_1 _4693_ (.A0(_2291_),
    .A1(_2292_),
    .S(net372),
    .X(_2293_));
 sky130_fd_sc_hd__mux4_1 _4694_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net391),
    .S1(net380),
    .X(_2294_));
 sky130_fd_sc_hd__mux4_1 _4695_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net390),
    .S1(net379),
    .X(_2295_));
 sky130_fd_sc_hd__mux2_1 _4696_ (.A0(_2295_),
    .A1(_2294_),
    .S(net372),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(_2296_),
    .A1(_2293_),
    .S(net368),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_1 _4698_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net389),
    .S1(net376),
    .X(_2297_));
 sky130_fd_sc_hd__mux4_1 _4699_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net389),
    .S1(net378),
    .X(_2298_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(_2297_),
    .A1(_2298_),
    .S(net371),
    .X(_2299_));
 sky130_fd_sc_hd__mux4_1 _4701_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net389),
    .S1(net376),
    .X(_2300_));
 sky130_fd_sc_hd__mux4_1 _4702_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net389),
    .S1(net376),
    .X(_2301_));
 sky130_fd_sc_hd__mux2_1 _4703_ (.A0(_2301_),
    .A1(_2300_),
    .S(net371),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_1 _4704_ (.A0(_2302_),
    .A1(_2299_),
    .S(net368),
    .X(_0002_));
 sky130_fd_sc_hd__mux4_1 _4705_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net396),
    .S1(net383),
    .X(_2303_));
 sky130_fd_sc_hd__mux4_1 _4706_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net396),
    .S1(net383),
    .X(_2304_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(_2303_),
    .A1(_2304_),
    .S(net374),
    .X(_2305_));
 sky130_fd_sc_hd__mux4_1 _4708_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net396),
    .S1(net383),
    .X(_2306_));
 sky130_fd_sc_hd__mux4_1 _4709_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net396),
    .S1(net383),
    .X(_2307_));
 sky130_fd_sc_hd__mux2_1 _4710_ (.A0(_2307_),
    .A1(_2306_),
    .S(net374),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(_2308_),
    .A1(_2305_),
    .S(net369),
    .X(_0003_));
 sky130_fd_sc_hd__mux4_1 _4712_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net390),
    .S1(net379),
    .X(_2309_));
 sky130_fd_sc_hd__mux4_1 _4713_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net390),
    .S1(net379),
    .X(_2310_));
 sky130_fd_sc_hd__mux2_1 _4714_ (.A0(_2309_),
    .A1(_2310_),
    .S(net372),
    .X(_2311_));
 sky130_fd_sc_hd__mux4_1 _4715_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net390),
    .S1(net379),
    .X(_2312_));
 sky130_fd_sc_hd__mux4_1 _4716_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net390),
    .S1(net379),
    .X(_2313_));
 sky130_fd_sc_hd__mux2_1 _4717_ (.A0(_2313_),
    .A1(_2312_),
    .S(net372),
    .X(_2314_));
 sky130_fd_sc_hd__mux2_1 _4718_ (.A0(_2314_),
    .A1(_2311_),
    .S(net368),
    .X(_0004_));
 sky130_fd_sc_hd__mux4_1 _4719_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net396),
    .S1(net385),
    .X(_2315_));
 sky130_fd_sc_hd__mux4_1 _4720_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net396),
    .S1(net385),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(_2315_),
    .A1(_2316_),
    .S(net374),
    .X(_2317_));
 sky130_fd_sc_hd__mux4_1 _4722_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net396),
    .S1(net385),
    .X(_2318_));
 sky130_fd_sc_hd__mux4_1 _4723_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net396),
    .S1(net385),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_1 _4724_ (.A0(_2319_),
    .A1(_2318_),
    .S(net374),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_1 _4725_ (.A0(_2320_),
    .A1(_2317_),
    .S(net369),
    .X(_0005_));
 sky130_fd_sc_hd__mux4_1 _4726_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net397),
    .S1(net382),
    .X(_2321_));
 sky130_fd_sc_hd__mux4_1 _4727_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net397),
    .S1(net382),
    .X(_2322_));
 sky130_fd_sc_hd__mux2_1 _4728_ (.A0(_2321_),
    .A1(_2322_),
    .S(net373),
    .X(_2323_));
 sky130_fd_sc_hd__mux4_1 _4729_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net396),
    .S1(net385),
    .X(_2324_));
 sky130_fd_sc_hd__mux4_1 _4730_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net397),
    .S1(net382),
    .X(_2325_));
 sky130_fd_sc_hd__mux2_1 _4731_ (.A0(_2325_),
    .A1(_2324_),
    .S(net373),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _4732_ (.A0(_2326_),
    .A1(_2323_),
    .S(net369),
    .X(_0006_));
 sky130_fd_sc_hd__mux4_1 _4733_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net391),
    .S1(net380),
    .X(_2327_));
 sky130_fd_sc_hd__mux4_1 _4734_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net392),
    .S1(net381),
    .X(_2328_));
 sky130_fd_sc_hd__mux2_1 _4735_ (.A0(_2327_),
    .A1(_2328_),
    .S(net373),
    .X(_2329_));
 sky130_fd_sc_hd__mux4_1 _4736_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net390),
    .S1(net380),
    .X(_2330_));
 sky130_fd_sc_hd__mux4_1 _4737_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net392),
    .S1(net381),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(_2331_),
    .A1(_2330_),
    .S(net373),
    .X(_2332_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(_2332_),
    .A1(_2329_),
    .S(net369),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _4740_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net393),
    .S1(net382),
    .X(_2333_));
 sky130_fd_sc_hd__mux4_1 _4741_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net393),
    .S1(net382),
    .X(_2334_));
 sky130_fd_sc_hd__mux2_1 _4742_ (.A0(_2333_),
    .A1(_2334_),
    .S(net373),
    .X(_2335_));
 sky130_fd_sc_hd__mux4_1 _4743_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net392),
    .S1(net382),
    .X(_2336_));
 sky130_fd_sc_hd__mux4_1 _4744_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net392),
    .S1(net382),
    .X(_2337_));
 sky130_fd_sc_hd__mux2_1 _4745_ (.A0(_2337_),
    .A1(_2336_),
    .S(net373),
    .X(_2338_));
 sky130_fd_sc_hd__mux2_1 _4746_ (.A0(_2338_),
    .A1(_2335_),
    .S(net369),
    .X(_0008_));
 sky130_fd_sc_hd__mux4_1 _4747_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net394),
    .S1(net383),
    .X(_2339_));
 sky130_fd_sc_hd__mux4_1 _4748_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net394),
    .S1(net383),
    .X(_2340_));
 sky130_fd_sc_hd__mux2_1 _4749_ (.A0(_2339_),
    .A1(_2340_),
    .S(net374),
    .X(_2341_));
 sky130_fd_sc_hd__mux4_1 _4750_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net394),
    .S1(net383),
    .X(_2342_));
 sky130_fd_sc_hd__mux4_1 _4751_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net394),
    .S1(net383),
    .X(_2343_));
 sky130_fd_sc_hd__mux2_1 _4752_ (.A0(_2343_),
    .A1(_2342_),
    .S(net374),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _4753_ (.A0(_2344_),
    .A1(_2341_),
    .S(net370),
    .X(_0009_));
 sky130_fd_sc_hd__mux4_1 _4754_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net390),
    .S1(net379),
    .X(_2345_));
 sky130_fd_sc_hd__mux4_1 _4755_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net390),
    .S1(net379),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(_2345_),
    .A1(_2346_),
    .S(net372),
    .X(_2347_));
 sky130_fd_sc_hd__mux4_1 _4757_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net390),
    .S1(net379),
    .X(_2348_));
 sky130_fd_sc_hd__mux4_1 _4758_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net390),
    .S1(net379),
    .X(_2349_));
 sky130_fd_sc_hd__mux2_1 _4759_ (.A0(_2349_),
    .A1(_2348_),
    .S(net372),
    .X(_2350_));
 sky130_fd_sc_hd__mux2_1 _4760_ (.A0(_2350_),
    .A1(_2347_),
    .S(net370),
    .X(_0010_));
 sky130_fd_sc_hd__mux4_1 _4761_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net388),
    .S1(net378),
    .X(_2351_));
 sky130_fd_sc_hd__mux4_1 _4762_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net388),
    .S1(net378),
    .X(_2352_));
 sky130_fd_sc_hd__mux2_1 _4763_ (.A0(_2351_),
    .A1(_2352_),
    .S(net371),
    .X(_2353_));
 sky130_fd_sc_hd__mux4_1 _4764_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net388),
    .S1(net386),
    .X(_2354_));
 sky130_fd_sc_hd__mux4_1 _4765_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net388),
    .S1(net386),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(_2355_),
    .A1(_2354_),
    .S(net371),
    .X(_2356_));
 sky130_fd_sc_hd__mux2_1 _4767_ (.A0(_2356_),
    .A1(_2353_),
    .S(net368),
    .X(_0012_));
 sky130_fd_sc_hd__mux4_1 _4768_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net388),
    .S1(net378),
    .X(_2357_));
 sky130_fd_sc_hd__mux4_1 _4769_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net388),
    .S1(net378),
    .X(_2358_));
 sky130_fd_sc_hd__mux2_1 _4770_ (.A0(_2357_),
    .A1(_2358_),
    .S(net371),
    .X(_2359_));
 sky130_fd_sc_hd__mux4_1 _4771_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net388),
    .S1(net378),
    .X(_2360_));
 sky130_fd_sc_hd__mux4_1 _4772_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net388),
    .S1(net378),
    .X(_2361_));
 sky130_fd_sc_hd__mux2_1 _4773_ (.A0(_2361_),
    .A1(_2360_),
    .S(net372),
    .X(_2362_));
 sky130_fd_sc_hd__mux2_1 _4774_ (.A0(_2362_),
    .A1(_2359_),
    .S(net368),
    .X(_0013_));
 sky130_fd_sc_hd__mux4_1 _4775_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net392),
    .S1(net381),
    .X(_2363_));
 sky130_fd_sc_hd__mux4_1 _4776_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net392),
    .S1(net381),
    .X(_2364_));
 sky130_fd_sc_hd__mux2_1 _4777_ (.A0(_2363_),
    .A1(_2364_),
    .S(net373),
    .X(_2365_));
 sky130_fd_sc_hd__mux4_1 _4778_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net392),
    .S1(net381),
    .X(_2366_));
 sky130_fd_sc_hd__mux4_1 _4779_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net392),
    .S1(net381),
    .X(_2367_));
 sky130_fd_sc_hd__mux2_1 _4780_ (.A0(_2367_),
    .A1(_2366_),
    .S(net373),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _4781_ (.A0(_2368_),
    .A1(_2365_),
    .S(net369),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_1 _4782_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net387),
    .S1(net376),
    .X(_2369_));
 sky130_fd_sc_hd__mux4_1 _4783_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net387),
    .S1(net376),
    .X(_2370_));
 sky130_fd_sc_hd__mux2_1 _4784_ (.A0(_2369_),
    .A1(_2370_),
    .S(net371),
    .X(_2371_));
 sky130_fd_sc_hd__mux4_1 _4785_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net387),
    .S1(net377),
    .X(_2372_));
 sky130_fd_sc_hd__mux4_1 _4786_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net387),
    .S1(net377),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_1 _4787_ (.A0(_2373_),
    .A1(_2372_),
    .S(net371),
    .X(_2374_));
 sky130_fd_sc_hd__mux2_1 _4788_ (.A0(_2374_),
    .A1(_2371_),
    .S(net368),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_1 _4789_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net394),
    .S1(net384),
    .X(_2375_));
 sky130_fd_sc_hd__mux4_1 _4790_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net394),
    .S1(net384),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_1 _4791_ (.A0(_2375_),
    .A1(_2376_),
    .S(net374),
    .X(_2377_));
 sky130_fd_sc_hd__mux4_1 _4792_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net394),
    .S1(net383),
    .X(_2378_));
 sky130_fd_sc_hd__mux4_1 _4793_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net394),
    .S1(net384),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_1 _4794_ (.A0(_2379_),
    .A1(_2378_),
    .S(net374),
    .X(_2380_));
 sky130_fd_sc_hd__mux2_1 _4795_ (.A0(_2380_),
    .A1(_2377_),
    .S(net370),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_1 _4796_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net387),
    .S1(net376),
    .X(_2381_));
 sky130_fd_sc_hd__mux4_1 _4797_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net387),
    .S1(net377),
    .X(_2382_));
 sky130_fd_sc_hd__mux2_1 _4798_ (.A0(_2381_),
    .A1(_2382_),
    .S(net371),
    .X(_2383_));
 sky130_fd_sc_hd__mux4_1 _4799_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net387),
    .S1(net377),
    .X(_2384_));
 sky130_fd_sc_hd__mux4_1 _4800_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net387),
    .S1(net377),
    .X(_2385_));
 sky130_fd_sc_hd__mux2_1 _4801_ (.A0(_2385_),
    .A1(_2384_),
    .S(net371),
    .X(_2386_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(_2386_),
    .A1(_2383_),
    .S(net368),
    .X(_0017_));
 sky130_fd_sc_hd__mux4_1 _4803_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net387),
    .S1(net377),
    .X(_2387_));
 sky130_fd_sc_hd__mux4_1 _4804_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net387),
    .S1(net377),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_1 _4805_ (.A0(_2387_),
    .A1(_2388_),
    .S(net371),
    .X(_2389_));
 sky130_fd_sc_hd__mux4_1 _4806_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net388),
    .S1(net377),
    .X(_2390_));
 sky130_fd_sc_hd__mux4_1 _4807_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net387),
    .S1(net377),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _4808_ (.A0(_2391_),
    .A1(_2390_),
    .S(net371),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _4809_ (.A0(_2392_),
    .A1(_2389_),
    .S(net368),
    .X(_0018_));
 sky130_fd_sc_hd__mux4_1 _4810_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net391),
    .S1(net379),
    .X(_2393_));
 sky130_fd_sc_hd__mux4_1 _4811_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net391),
    .S1(net379),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(_2393_),
    .A1(_2394_),
    .S(net372),
    .X(_2395_));
 sky130_fd_sc_hd__mux4_1 _4813_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net391),
    .S1(net380),
    .X(_2396_));
 sky130_fd_sc_hd__mux4_1 _4814_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net391),
    .S1(net380),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _4815_ (.A0(_2397_),
    .A1(_2396_),
    .S(net372),
    .X(_2398_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(_2398_),
    .A1(_2395_),
    .S(net368),
    .X(_0019_));
 sky130_fd_sc_hd__mux4_1 _4817_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net389),
    .S1(net376),
    .X(_2399_));
 sky130_fd_sc_hd__mux4_1 _4818_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net389),
    .S1(net376),
    .X(_2400_));
 sky130_fd_sc_hd__mux2_1 _4819_ (.A0(_2399_),
    .A1(_2400_),
    .S(net371),
    .X(_2401_));
 sky130_fd_sc_hd__mux4_1 _4820_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net389),
    .S1(net376),
    .X(_2402_));
 sky130_fd_sc_hd__mux4_1 _4821_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net389),
    .S1(net376),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_2403_),
    .A1(_2402_),
    .S(net371),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(_2404_),
    .A1(_2401_),
    .S(net368),
    .X(_0020_));
 sky130_fd_sc_hd__mux4_1 _4824_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net387),
    .S1(net376),
    .X(_2405_));
 sky130_fd_sc_hd__mux4_1 _4825_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net387),
    .S1(net376),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_1 _4826_ (.A0(_2405_),
    .A1(_2406_),
    .S(net371),
    .X(_2407_));
 sky130_fd_sc_hd__mux4_1 _4827_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net387),
    .S1(net376),
    .X(_2408_));
 sky130_fd_sc_hd__mux4_1 _4828_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net387),
    .S1(net376),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _4829_ (.A0(_2409_),
    .A1(_2408_),
    .S(net371),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _4830_ (.A0(_2410_),
    .A1(_2407_),
    .S(net368),
    .X(_0021_));
 sky130_fd_sc_hd__mux4_1 _4831_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net388),
    .S1(net378),
    .X(_2411_));
 sky130_fd_sc_hd__mux4_1 _4832_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net388),
    .S1(net378),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _4833_ (.A0(_2411_),
    .A1(_2412_),
    .S(net372),
    .X(_2413_));
 sky130_fd_sc_hd__mux4_1 _4834_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net388),
    .S1(net378),
    .X(_2414_));
 sky130_fd_sc_hd__mux4_1 _4835_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net390),
    .S1(net379),
    .X(_2415_));
 sky130_fd_sc_hd__mux2_1 _4836_ (.A0(_2415_),
    .A1(_2414_),
    .S(net372),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _4837_ (.A0(_2416_),
    .A1(_2413_),
    .S(net368),
    .X(_0023_));
 sky130_fd_sc_hd__mux4_1 _4838_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net388),
    .S1(net378),
    .X(_2417_));
 sky130_fd_sc_hd__mux4_1 _4839_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net388),
    .S1(net378),
    .X(_2418_));
 sky130_fd_sc_hd__mux2_1 _4840_ (.A0(_2417_),
    .A1(_2418_),
    .S(net372),
    .X(_2419_));
 sky130_fd_sc_hd__mux4_1 _4841_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net388),
    .S1(net378),
    .X(_2420_));
 sky130_fd_sc_hd__mux4_1 _4842_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net387),
    .S1(net376),
    .X(_2421_));
 sky130_fd_sc_hd__mux2_1 _4843_ (.A0(_2421_),
    .A1(_2420_),
    .S(net372),
    .X(_2422_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(_2422_),
    .A1(_2419_),
    .S(net368),
    .X(_0024_));
 sky130_fd_sc_hd__and3_1 _4845_ (.A(_1301_),
    .B(net248),
    .C(net2131),
    .X(_2423_));
 sky130_fd_sc_hd__nand2_1 _4846_ (.A(net249),
    .B(net183),
    .Y(_2424_));
 sky130_fd_sc_hd__nor2_1 _4847_ (.A(_1277_),
    .B(net163),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_2 _4848_ (.A(net578),
    .B(net2038),
    .Y(_2425_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(net2018),
    .B(net920),
    .Y(_2426_));
 sky130_fd_sc_hd__a21oi_1 _4850_ (.A1(net579),
    .A2(net2019),
    .B1(net163),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _4851_ (.A(net2106),
    .B(net920),
    .Y(_2427_));
 sky130_fd_sc_hd__a21oi_4 _4852_ (.A1(_2425_),
    .A2(_2427_),
    .B1(net162),
    .Y(_0195_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(net1924),
    .B(net920),
    .Y(_2428_));
 sky130_fd_sc_hd__a21oi_1 _4854_ (.A1(net579),
    .A2(net1925),
    .B1(net163),
    .Y(_0196_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(net587),
    .B(_2036_),
    .Y(_2429_));
 sky130_fd_sc_hd__a21oi_1 _4856_ (.A1(net579),
    .A2(net588),
    .B1(net162),
    .Y(_0197_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(net2056),
    .B(net920),
    .Y(_2430_));
 sky130_fd_sc_hd__a21oi_1 _4858_ (.A1(net579),
    .A2(net2057),
    .B1(net163),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _4859_ (.A(net708),
    .B(net920),
    .Y(_2431_));
 sky130_fd_sc_hd__a21oi_1 _4860_ (.A1(net579),
    .A2(_2431_),
    .B1(net163),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(net2221),
    .B(_2036_),
    .Y(_2432_));
 sky130_fd_sc_hd__a21oi_1 _4862_ (.A1(net579),
    .A2(_2432_),
    .B1(net162),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(net368),
    .B(net920),
    .Y(_2433_));
 sky130_fd_sc_hd__a21oi_1 _4864_ (.A1(net579),
    .A2(net1190),
    .B1(net163),
    .Y(_0201_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(net371),
    .B(net920),
    .Y(_2434_));
 sky130_fd_sc_hd__a21oi_1 _4866_ (.A1(net579),
    .A2(net2055),
    .B1(net163),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(net376),
    .B(net920),
    .Y(_2435_));
 sky130_fd_sc_hd__a21oi_1 _4868_ (.A1(net579),
    .A2(net921),
    .B1(net163),
    .Y(_0203_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(net389),
    .B(net920),
    .Y(_2436_));
 sky130_fd_sc_hd__a21oi_1 _4870_ (.A1(net579),
    .A2(net1715),
    .B1(net163),
    .Y(_0204_));
 sky130_fd_sc_hd__a21o_4 _4871_ (.A1(net2037),
    .A2(_2034_),
    .B1(net920),
    .X(_2437_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(net2020),
    .B(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__or2_4 _4873_ (.A(_1277_),
    .B(_2437_),
    .X(_2439_));
 sky130_fd_sc_hd__a21oi_1 _4874_ (.A1(net2021),
    .A2(_2439_),
    .B1(net162),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_1 _4875_ (.A(net398),
    .B(_2437_),
    .Y(_2440_));
 sky130_fd_sc_hd__a21oi_1 _4876_ (.A1(_2439_),
    .A2(_2440_),
    .B1(net162),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _4877_ (.A(net2234),
    .B(_2437_),
    .Y(_2441_));
 sky130_fd_sc_hd__a21oi_1 _4878_ (.A1(_2439_),
    .A2(_2441_),
    .B1(net162),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(net410),
    .B(_2437_),
    .Y(_2442_));
 sky130_fd_sc_hd__a21oi_1 _4880_ (.A1(_2439_),
    .A2(_2442_),
    .B1(net162),
    .Y(_0208_));
 sky130_fd_sc_hd__nand2_1 _4881_ (.A(net422),
    .B(_2437_),
    .Y(_2443_));
 sky130_fd_sc_hd__a21oi_1 _4882_ (.A1(_2439_),
    .A2(_2443_),
    .B1(net162),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(net2119),
    .B(_2437_),
    .Y(_2444_));
 sky130_fd_sc_hd__a21oi_1 _4884_ (.A1(_2439_),
    .A2(_2444_),
    .B1(net162),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(net2148),
    .B(_2437_),
    .Y(_2445_));
 sky130_fd_sc_hd__a21oi_1 _4886_ (.A1(_2439_),
    .A2(_2445_),
    .B1(net163),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(net2095),
    .B(_2437_),
    .Y(_2446_));
 sky130_fd_sc_hd__a21oi_1 _4888_ (.A1(_2439_),
    .A2(_2446_),
    .B1(net162),
    .Y(_0212_));
 sky130_fd_sc_hd__and3b_4 _4889_ (.A_N(net919),
    .B(_2032_),
    .C(net2029),
    .X(_2447_));
 sky130_fd_sc_hd__and2_1 _4890_ (.A(_1280_),
    .B(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__nor2_1 _4891_ (.A(_2437_),
    .B(_2447_),
    .Y(_2449_));
 sky130_fd_sc_hd__o21a_1 _4892_ (.A1(_2448_),
    .A2(_2449_),
    .B1(net578),
    .X(_2450_));
 sky130_fd_sc_hd__and3_1 _4893_ (.A(net397),
    .B(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ),
    .C(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .X(_2451_));
 sky130_fd_sc_hd__a21o_1 _4894_ (.A1(net1959),
    .A2(_2032_),
    .B1(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__and4b_1 _4895_ (.A_N(net919),
    .B(_2452_),
    .C(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .D(net2029),
    .X(_2453_));
 sky130_fd_sc_hd__o21a_1 _4896_ (.A1(_2450_),
    .A2(net2030),
    .B1(net176),
    .X(_0213_));
 sky130_fd_sc_hd__and3_1 _4897_ (.A(net2018),
    .B(net2038),
    .C(net176),
    .X(_0214_));
 sky130_fd_sc_hd__and3_1 _4898_ (.A(net2106),
    .B(net2038),
    .C(net175),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _4899_ (.A(net1924),
    .B(net2038),
    .C(net176),
    .X(_0216_));
 sky130_fd_sc_hd__and3_1 _4900_ (.A(net587),
    .B(net2038),
    .C(net175),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _4901_ (.A(net2056),
    .B(net2038),
    .C(net175),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _4902_ (.A(net708),
    .B(_2037_),
    .C(net175),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_2 _4903_ (.A1(net2037),
    .A2(_2034_),
    .B1(_2449_),
    .X(_2454_));
 sky130_fd_sc_hd__a22o_1 _4904_ (.A1(net2127),
    .A2(_2447_),
    .B1(_2454_),
    .B2(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ),
    .X(_2455_));
 sky130_fd_sc_hd__and2_1 _4905_ (.A(net175),
    .B(net2128),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _4906_ (.A1(net608),
    .A2(_2447_),
    .B1(_2454_),
    .B2(net369),
    .X(_2456_));
 sky130_fd_sc_hd__and2_1 _4907_ (.A(net176),
    .B(_2456_),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_1 _4908_ (.A1(net2042),
    .A2(_2447_),
    .B1(_2454_),
    .B2(net373),
    .X(_2457_));
 sky130_fd_sc_hd__and2_1 _4909_ (.A(net175),
    .B(_2457_),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _4910_ (.A1(net1946),
    .A2(_2447_),
    .B1(_2454_),
    .B2(net381),
    .X(_2458_));
 sky130_fd_sc_hd__and2_1 _4911_ (.A(net175),
    .B(_2458_),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _4912_ (.A1(net1959),
    .A2(_2448_),
    .B1(_2449_),
    .B2(net397),
    .X(_2459_));
 sky130_fd_sc_hd__and2_1 _4913_ (.A(net176),
    .B(_2459_),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_1 _4914_ (.A(net2148),
    .B(net426),
    .Y(_2460_));
 sky130_fd_sc_hd__nand2_2 _4915_ (.A(_1278_),
    .B(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__and3_1 _4916_ (.A(_1280_),
    .B(_1281_),
    .C(_2032_),
    .X(_2462_));
 sky130_fd_sc_hd__o2111ai_4 _4917_ (.A1(_1281_),
    .A2(_2461_),
    .B1(net919),
    .C1(_1280_),
    .D1(_2032_),
    .Y(_2463_));
 sky130_fd_sc_hd__inv_2 _4918_ (.A(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__or4_4 _4919_ (.A(_2038_),
    .B(_2447_),
    .C(_2462_),
    .D(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__or3_1 _4920_ (.A(net2018),
    .B(_2461_),
    .C(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__o21a_1 _4921_ (.A1(_2461_),
    .A2(_2463_),
    .B1(_2465_),
    .X(_2467_));
 sky130_fd_sc_hd__or4b_1 _4922_ (.A(net2119),
    .B(net2148),
    .C(_2463_),
    .D_N(net426),
    .X(_2468_));
 sky130_fd_sc_hd__or4_1 _4923_ (.A(net2119),
    .B(_1279_),
    .C(net426),
    .D(_2463_),
    .X(_2469_));
 sky130_fd_sc_hd__or4b_2 _4924_ (.A(_1278_),
    .B(net2148),
    .C(_2463_),
    .D_N(net426),
    .X(_2470_));
 sky130_fd_sc_hd__and4_1 _4925_ (.A(net2287),
    .B(net2248),
    .C(net426),
    .D(_2464_),
    .X(_2471_));
 sky130_fd_sc_hd__or4_1 _4926_ (.A(_1278_),
    .B(_1279_),
    .C(net426),
    .D(_2463_),
    .X(_2472_));
 sky130_fd_sc_hd__o211a_1 _4927_ (.A1(net2248),
    .A2(net426),
    .B1(_2464_),
    .C1(net2119),
    .X(_2473_));
 sky130_fd_sc_hd__nand2_2 _4928_ (.A(net2029),
    .B(_2036_),
    .Y(_2474_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__and2_1 _4930_ (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .B(_2447_),
    .X(_2476_));
 sky130_fd_sc_hd__nand2_2 _4931_ (.A(net2170),
    .B(_2447_),
    .Y(_2477_));
 sky130_fd_sc_hd__and4_1 _4932_ (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .B(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .C(net426),
    .D(_2476_),
    .X(_2478_));
 sky130_fd_sc_hd__or4_1 _4933_ (.A(_1278_),
    .B(_1279_),
    .C(net426),
    .D(_2477_),
    .X(_2479_));
 sky130_fd_sc_hd__or3_1 _4934_ (.A(_1278_),
    .B(net426),
    .C(_2477_),
    .X(_2480_));
 sky130_fd_sc_hd__o2bb2a_1 _4935_ (.A1_N(_0066_),
    .A2_N(_2474_),
    .B1(_2477_),
    .B2(_1278_),
    .X(_2481_));
 sky130_fd_sc_hd__or4b_1 _4936_ (.A(net2287),
    .B(_2477_),
    .C(net2286),
    .D_N(net426),
    .X(_2482_));
 sky130_fd_sc_hd__and3_1 _4937_ (.A(_1278_),
    .B(_1279_),
    .C(_2476_),
    .X(_2483_));
 sky130_fd_sc_hd__o32a_1 _4938_ (.A1(_2473_),
    .A2(_2481_),
    .A3(_2483_),
    .B1(_2470_),
    .B2(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ),
    .X(_2484_));
 sky130_fd_sc_hd__or3b_1 _4939_ (.A(_1278_),
    .B(_2463_),
    .C_N(_2460_),
    .X(_2485_));
 sky130_fd_sc_hd__inv_2 _4940_ (.A(_2485_),
    .Y(_2486_));
 sky130_fd_sc_hd__and4_1 _4941_ (.A(_1278_),
    .B(net2148),
    .C(net426),
    .D(_2464_),
    .X(_2487_));
 sky130_fd_sc_hd__o311a_1 _4942_ (.A1(_2484_),
    .A2(_2486_),
    .A3(_2487_),
    .B1(_2469_),
    .C1(_2468_),
    .X(_2488_));
 sky130_fd_sc_hd__inv_2 _4943_ (.A(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__a2bb2o_1 _4944_ (.A1_N(_2461_),
    .A2_N(_2465_),
    .B1(_2467_),
    .B2(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__and3_1 _4945_ (.A(net174),
    .B(_2466_),
    .C(_2490_),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _4946_ (.A(_2467_),
    .B(_2468_),
    .C(_2469_),
    .X(_2491_));
 sky130_fd_sc_hd__a21oi_1 _4947_ (.A1(_0064_),
    .A2(_2474_),
    .B1(_2478_),
    .Y(_2492_));
 sky130_fd_sc_hd__a41o_1 _4948_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .A2(_1279_),
    .A3(net426),
    .A4(_2476_),
    .B1(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__a32o_1 _4949_ (.A1(net2288),
    .A2(_2460_),
    .A3(_2476_),
    .B1(_2479_),
    .B2(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__a2bb2o_1 _4950_ (.A1_N(_2461_),
    .A2_N(_2477_),
    .B1(_2482_),
    .B2(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__o211a_1 _4951_ (.A1(_2471_),
    .A2(_2495_),
    .B1(_2472_),
    .C1(_2470_),
    .X(_2496_));
 sky130_fd_sc_hd__o21a_1 _4952_ (.A1(net2018),
    .A2(_2470_),
    .B1(_2485_),
    .X(_2497_));
 sky130_fd_sc_hd__or3b_1 _4953_ (.A(_2487_),
    .B(_2496_),
    .C_N(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a2bb2o_1 _4954_ (.A1_N(_2461_),
    .A2_N(_2465_),
    .B1(_2491_),
    .B2(_2498_),
    .X(_2499_));
 sky130_fd_sc_hd__a21oi_1 _4955_ (.A1(_2466_),
    .A2(_2499_),
    .B1(net162),
    .Y(_0226_));
 sky130_fd_sc_hd__a32o_1 _4956_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .A2(net426),
    .A3(_2476_),
    .B1(_2474_),
    .B2(_0065_),
    .X(_2500_));
 sky130_fd_sc_hd__a21oi_1 _4957_ (.A1(_2480_),
    .A2(_2500_),
    .B1(_2483_),
    .Y(_2501_));
 sky130_fd_sc_hd__o21a_1 _4958_ (.A1(_2473_),
    .A2(_2501_),
    .B1(_2497_),
    .X(_2502_));
 sky130_fd_sc_hd__o21ai_1 _4959_ (.A1(_2487_),
    .A2(_2502_),
    .B1(_2469_),
    .Y(_2503_));
 sky130_fd_sc_hd__nand2_1 _4960_ (.A(_2468_),
    .B(_2503_),
    .Y(_2504_));
 sky130_fd_sc_hd__a2bb2o_1 _4961_ (.A1_N(_2461_),
    .A2_N(_2465_),
    .B1(_2467_),
    .B2(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__a21oi_1 _4962_ (.A1(_2466_),
    .A2(_2505_),
    .B1(net162),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _4963_ (.A(_2033_),
    .B(net2038),
    .Y(_2506_));
 sky130_fd_sc_hd__and3_1 _4964_ (.A(_1281_),
    .B(net175),
    .C(_2506_),
    .X(_0228_));
 sky130_fd_sc_hd__or2_4 _4965_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_2507_));
 sky130_fd_sc_hd__nor2_1 _4966_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_2508_));
 sky130_fd_sc_hd__or4bb_4 _4967_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(net464),
    .C_N(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .D_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .X(_2509_));
 sky130_fd_sc_hd__nor2_4 _4968_ (.A(_2507_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__or2_4 _4969_ (.A(_2507_),
    .B(_2509_),
    .X(_2511_));
 sky130_fd_sc_hd__or3_1 _4970_ (.A(net464),
    .B(net2096),
    .C(net330),
    .X(_2512_));
 sky130_fd_sc_hd__o21a_1 _4971_ (.A1(net298),
    .A2(net327),
    .B1(_2512_),
    .X(_0229_));
 sky130_fd_sc_hd__and2_1 _4972_ (.A(net299),
    .B(net330),
    .X(_2513_));
 sky130_fd_sc_hd__a31o_1 _4973_ (.A1(net447),
    .A2(net1836),
    .A3(net327),
    .B1(_2513_),
    .X(_0230_));
 sky130_fd_sc_hd__and2_1 _4974_ (.A(net353),
    .B(net330),
    .X(_2514_));
 sky130_fd_sc_hd__a31o_1 _4975_ (.A1(net447),
    .A2(net1882),
    .A3(net327),
    .B1(_2514_),
    .X(_0231_));
 sky130_fd_sc_hd__and2_1 _4976_ (.A(net355),
    .B(net330),
    .X(_2515_));
 sky130_fd_sc_hd__a31o_1 _4977_ (.A1(net454),
    .A2(net1902),
    .A3(net327),
    .B1(_2515_),
    .X(_0232_));
 sky130_fd_sc_hd__and2_1 _4978_ (.A(net356),
    .B(net330),
    .X(_2516_));
 sky130_fd_sc_hd__a31o_1 _4979_ (.A1(net452),
    .A2(net1832),
    .A3(net327),
    .B1(_2516_),
    .X(_0233_));
 sky130_fd_sc_hd__and2_1 _4980_ (.A(net354),
    .B(net330),
    .X(_2517_));
 sky130_fd_sc_hd__a31o_1 _4981_ (.A1(net452),
    .A2(net1805),
    .A3(net327),
    .B1(_2517_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _4982_ (.A(net352),
    .B(net329),
    .X(_2518_));
 sky130_fd_sc_hd__a31o_1 _4983_ (.A1(net439),
    .A2(net1645),
    .A3(net328),
    .B1(_2518_),
    .X(_0235_));
 sky130_fd_sc_hd__and2_1 _4984_ (.A(net351),
    .B(net330),
    .X(_2519_));
 sky130_fd_sc_hd__a31o_1 _4985_ (.A1(net445),
    .A2(net1838),
    .A3(net327),
    .B1(_2519_),
    .X(_0236_));
 sky130_fd_sc_hd__and2_1 _4986_ (.A(net358),
    .B(net329),
    .X(_2520_));
 sky130_fd_sc_hd__a31o_1 _4987_ (.A1(net446),
    .A2(net1876),
    .A3(net328),
    .B1(_2520_),
    .X(_0237_));
 sky130_fd_sc_hd__and2_1 _4988_ (.A(net359),
    .B(net330),
    .X(_2521_));
 sky130_fd_sc_hd__a31o_1 _4989_ (.A1(net456),
    .A2(net1746),
    .A3(net327),
    .B1(_2521_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_1 _4990_ (.A(net357),
    .B(net329),
    .X(_2522_));
 sky130_fd_sc_hd__a31o_1 _4991_ (.A1(net439),
    .A2(net2001),
    .A3(net328),
    .B1(_2522_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _4992_ (.A(net361),
    .B(net329),
    .X(_2523_));
 sky130_fd_sc_hd__a31o_1 _4993_ (.A1(net430),
    .A2(net1763),
    .A3(net328),
    .B1(_2523_),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_1 _4994_ (.A(_1350_),
    .B(net327),
    .Y(_2524_));
 sky130_fd_sc_hd__a31o_1 _4995_ (.A1(net452),
    .A2(net1988),
    .A3(net327),
    .B1(_2524_),
    .X(_0241_));
 sky130_fd_sc_hd__and2_1 _4996_ (.A(net360),
    .B(net329),
    .X(_2525_));
 sky130_fd_sc_hd__a31o_1 _4997_ (.A1(net439),
    .A2(net1717),
    .A3(net328),
    .B1(_2525_),
    .X(_0242_));
 sky130_fd_sc_hd__and2_1 _4998_ (.A(net350),
    .B(net330),
    .X(_2526_));
 sky130_fd_sc_hd__a31o_1 _4999_ (.A1(net451),
    .A2(net1942),
    .A3(net327),
    .B1(_2526_),
    .X(_0243_));
 sky130_fd_sc_hd__and2_1 _5000_ (.A(net349),
    .B(net330),
    .X(_2527_));
 sky130_fd_sc_hd__a31o_1 _5001_ (.A1(net442),
    .A2(net1668),
    .A3(net327),
    .B1(_2527_),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _5002_ (.A(net345),
    .B(net330),
    .X(_2528_));
 sky130_fd_sc_hd__a31o_1 _5003_ (.A1(net445),
    .A2(net1759),
    .A3(net327),
    .B1(_2528_),
    .X(_0245_));
 sky130_fd_sc_hd__and2_1 _5004_ (.A(net344),
    .B(net330),
    .X(_2529_));
 sky130_fd_sc_hd__a31o_1 _5005_ (.A1(net448),
    .A2(net1787),
    .A3(net327),
    .B1(_2529_),
    .X(_0246_));
 sky130_fd_sc_hd__and2_1 _5006_ (.A(net341),
    .B(net330),
    .X(_2530_));
 sky130_fd_sc_hd__a31o_1 _5007_ (.A1(net455),
    .A2(net1870),
    .A3(_2511_),
    .B1(_2530_),
    .X(_0247_));
 sky130_fd_sc_hd__and2_1 _5008_ (.A(net343),
    .B(net329),
    .X(_2531_));
 sky130_fd_sc_hd__a31o_1 _5009_ (.A1(net438),
    .A2(net1934),
    .A3(net328),
    .B1(_2531_),
    .X(_0248_));
 sky130_fd_sc_hd__and2_1 _5010_ (.A(net342),
    .B(net329),
    .X(_2532_));
 sky130_fd_sc_hd__a31o_1 _5011_ (.A1(net433),
    .A2(net1765),
    .A3(net328),
    .B1(_2532_),
    .X(_0249_));
 sky130_fd_sc_hd__and2_1 _5012_ (.A(net346),
    .B(net329),
    .X(_2533_));
 sky130_fd_sc_hd__a31o_1 _5013_ (.A1(net437),
    .A2(net1816),
    .A3(net328),
    .B1(_2533_),
    .X(_0250_));
 sky130_fd_sc_hd__and2_1 _5014_ (.A(net348),
    .B(net330),
    .X(_2534_));
 sky130_fd_sc_hd__a31o_1 _5015_ (.A1(net445),
    .A2(net1752),
    .A3(net327),
    .B1(_2534_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_1 _5016_ (.A(net347),
    .B(net329),
    .X(_2535_));
 sky130_fd_sc_hd__a31o_1 _5017_ (.A1(net434),
    .A2(net1864),
    .A3(net328),
    .B1(_2535_),
    .X(_0252_));
 sky130_fd_sc_hd__and2_1 _5018_ (.A(net334),
    .B(net330),
    .X(_2536_));
 sky130_fd_sc_hd__a31o_1 _5019_ (.A1(net455),
    .A2(net1785),
    .A3(net327),
    .B1(_2536_),
    .X(_0253_));
 sky130_fd_sc_hd__and2_1 _5020_ (.A(net337),
    .B(net329),
    .X(_2537_));
 sky130_fd_sc_hd__a31o_1 _5021_ (.A1(net433),
    .A2(net1744),
    .A3(net328),
    .B1(_2537_),
    .X(_0254_));
 sky130_fd_sc_hd__and2_1 _5022_ (.A(net338),
    .B(net329),
    .X(_2538_));
 sky130_fd_sc_hd__a31o_1 _5023_ (.A1(net434),
    .A2(net1670),
    .A3(net328),
    .B1(_2538_),
    .X(_0255_));
 sky130_fd_sc_hd__and2_1 _5024_ (.A(net336),
    .B(net329),
    .X(_2539_));
 sky130_fd_sc_hd__a31o_1 _5025_ (.A1(net438),
    .A2(net1613),
    .A3(net328),
    .B1(_2539_),
    .X(_0256_));
 sky130_fd_sc_hd__and2_1 _5026_ (.A(net333),
    .B(net329),
    .X(_2540_));
 sky130_fd_sc_hd__a31o_1 _5027_ (.A1(net430),
    .A2(net1890),
    .A3(net328),
    .B1(_2540_),
    .X(_0257_));
 sky130_fd_sc_hd__and2_1 _5028_ (.A(net339),
    .B(net329),
    .X(_2541_));
 sky130_fd_sc_hd__a31o_1 _5029_ (.A1(net433),
    .A2(net1807),
    .A3(net328),
    .B1(_2541_),
    .X(_0258_));
 sky130_fd_sc_hd__and2_1 _5030_ (.A(net340),
    .B(net329),
    .X(_2542_));
 sky130_fd_sc_hd__a31o_1 _5031_ (.A1(net436),
    .A2(net1651),
    .A3(net328),
    .B1(_2542_),
    .X(_0259_));
 sky130_fd_sc_hd__and2_1 _5032_ (.A(net335),
    .B(net329),
    .X(_2543_));
 sky130_fd_sc_hd__a31o_1 _5033_ (.A1(net434),
    .A2(net1777),
    .A3(net328),
    .B1(_2543_),
    .X(_0260_));
 sky130_fd_sc_hd__or4b_4 _5034_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1286_),
    .C(net464),
    .D_N(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_2544_));
 sky130_fd_sc_hd__nor2_4 _5035_ (.A(_2507_),
    .B(_2544_),
    .Y(_2545_));
 sky130_fd_sc_hd__or2_4 _5036_ (.A(_2507_),
    .B(_2544_),
    .X(_2546_));
 sky130_fd_sc_hd__and2_1 _5037_ (.A(net298),
    .B(net297),
    .X(_2547_));
 sky130_fd_sc_hd__a31o_1 _5038_ (.A1(net454),
    .A2(net1769),
    .A3(net294),
    .B1(_2547_),
    .X(_0261_));
 sky130_fd_sc_hd__or3_1 _5039_ (.A(net464),
    .B(net2093),
    .C(net297),
    .X(_2548_));
 sky130_fd_sc_hd__o21a_1 _5040_ (.A1(net299),
    .A2(net294),
    .B1(_2548_),
    .X(_0262_));
 sky130_fd_sc_hd__and2_1 _5041_ (.A(net353),
    .B(net297),
    .X(_2549_));
 sky130_fd_sc_hd__a31o_1 _5042_ (.A1(net448),
    .A2(net1906),
    .A3(net294),
    .B1(_2549_),
    .X(_0263_));
 sky130_fd_sc_hd__and2_1 _5043_ (.A(net355),
    .B(net297),
    .X(_2550_));
 sky130_fd_sc_hd__a31o_1 _5044_ (.A1(net455),
    .A2(net1814),
    .A3(net294),
    .B1(_2550_),
    .X(_0264_));
 sky130_fd_sc_hd__and2_1 _5045_ (.A(net356),
    .B(net297),
    .X(_2551_));
 sky130_fd_sc_hd__a31o_1 _5046_ (.A1(net452),
    .A2(net1868),
    .A3(net294),
    .B1(_2551_),
    .X(_0265_));
 sky130_fd_sc_hd__and2_1 _5047_ (.A(net354),
    .B(net297),
    .X(_2552_));
 sky130_fd_sc_hd__a31o_1 _5048_ (.A1(net452),
    .A2(net1803),
    .A3(net294),
    .B1(_2552_),
    .X(_0266_));
 sky130_fd_sc_hd__and2_1 _5049_ (.A(net352),
    .B(net296),
    .X(_2553_));
 sky130_fd_sc_hd__a31o_1 _5050_ (.A1(net439),
    .A2(net1797),
    .A3(net295),
    .B1(_2553_),
    .X(_0267_));
 sky130_fd_sc_hd__and2_1 _5051_ (.A(net351),
    .B(net297),
    .X(_2554_));
 sky130_fd_sc_hd__a31o_1 _5052_ (.A1(net445),
    .A2(net1920),
    .A3(net294),
    .B1(_2554_),
    .X(_0268_));
 sky130_fd_sc_hd__and2_1 _5053_ (.A(net358),
    .B(net296),
    .X(_2555_));
 sky130_fd_sc_hd__a31o_1 _5054_ (.A1(net446),
    .A2(net1846),
    .A3(net295),
    .B1(_2555_),
    .X(_0269_));
 sky130_fd_sc_hd__and2_1 _5055_ (.A(net359),
    .B(net297),
    .X(_2556_));
 sky130_fd_sc_hd__a31o_1 _5056_ (.A1(net456),
    .A2(net1737),
    .A3(net294),
    .B1(_2556_),
    .X(_0270_));
 sky130_fd_sc_hd__and2_1 _5057_ (.A(net357),
    .B(net296),
    .X(_2557_));
 sky130_fd_sc_hd__a31o_1 _5058_ (.A1(net438),
    .A2(net1990),
    .A3(net295),
    .B1(_2557_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _5059_ (.A(net361),
    .B(net296),
    .X(_2558_));
 sky130_fd_sc_hd__a31o_1 _5060_ (.A1(net430),
    .A2(net1812),
    .A3(net295),
    .B1(_2558_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _5061_ (.A(_1350_),
    .B(_2546_),
    .Y(_2559_));
 sky130_fd_sc_hd__a31o_1 _5062_ (.A1(net452),
    .A2(net1848),
    .A3(net294),
    .B1(_2559_),
    .X(_0273_));
 sky130_fd_sc_hd__and2_1 _5063_ (.A(net360),
    .B(net296),
    .X(_2560_));
 sky130_fd_sc_hd__a31o_1 _5064_ (.A1(net439),
    .A2(net1896),
    .A3(net295),
    .B1(_2560_),
    .X(_0274_));
 sky130_fd_sc_hd__and2_1 _5065_ (.A(net350),
    .B(net297),
    .X(_2561_));
 sky130_fd_sc_hd__a31o_1 _5066_ (.A1(net451),
    .A2(net1912),
    .A3(net294),
    .B1(_2561_),
    .X(_0275_));
 sky130_fd_sc_hd__and2_1 _5067_ (.A(net349),
    .B(net297),
    .X(_2562_));
 sky130_fd_sc_hd__a31o_1 _5068_ (.A1(net443),
    .A2(net1842),
    .A3(net294),
    .B1(_2562_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _5069_ (.A(net345),
    .B(net297),
    .X(_2563_));
 sky130_fd_sc_hd__a31o_1 _5070_ (.A1(net445),
    .A2(net1880),
    .A3(net294),
    .B1(_2563_),
    .X(_0277_));
 sky130_fd_sc_hd__and2_1 _5071_ (.A(net344),
    .B(net297),
    .X(_2564_));
 sky130_fd_sc_hd__a31o_1 _5072_ (.A1(net448),
    .A2(net1854),
    .A3(net294),
    .B1(_2564_),
    .X(_0278_));
 sky130_fd_sc_hd__and2_1 _5073_ (.A(net341),
    .B(net297),
    .X(_2565_));
 sky130_fd_sc_hd__a31o_1 _5074_ (.A1(net455),
    .A2(net1826),
    .A3(net294),
    .B1(_2565_),
    .X(_0279_));
 sky130_fd_sc_hd__and2_1 _5075_ (.A(_1561_),
    .B(net296),
    .X(_2566_));
 sky130_fd_sc_hd__a31o_1 _5076_ (.A1(net438),
    .A2(net1904),
    .A3(net295),
    .B1(_2566_),
    .X(_0280_));
 sky130_fd_sc_hd__and2_1 _5077_ (.A(net342),
    .B(net296),
    .X(_2567_));
 sky130_fd_sc_hd__a31o_1 _5078_ (.A1(net436),
    .A2(net1773),
    .A3(net295),
    .B1(_2567_),
    .X(_0281_));
 sky130_fd_sc_hd__and2_1 _5079_ (.A(net346),
    .B(net296),
    .X(_2568_));
 sky130_fd_sc_hd__a31o_1 _5080_ (.A1(net437),
    .A2(net1820),
    .A3(net295),
    .B1(_2568_),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _5081_ (.A(net348),
    .B(net297),
    .X(_2569_));
 sky130_fd_sc_hd__a31o_1 _5082_ (.A1(net445),
    .A2(net1767),
    .A3(net294),
    .B1(_2569_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_1 _5083_ (.A(net347),
    .B(net296),
    .X(_2570_));
 sky130_fd_sc_hd__a31o_1 _5084_ (.A1(net433),
    .A2(net1754),
    .A3(net295),
    .B1(_2570_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _5085_ (.A(net334),
    .B(net297),
    .X(_2571_));
 sky130_fd_sc_hd__a31o_1 _5086_ (.A1(net455),
    .A2(net1872),
    .A3(net294),
    .B1(_2571_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_1 _5087_ (.A(net337),
    .B(net296),
    .X(_2572_));
 sky130_fd_sc_hd__a31o_1 _5088_ (.A1(net433),
    .A2(net1949),
    .A3(net295),
    .B1(_2572_),
    .X(_0286_));
 sky130_fd_sc_hd__and2_1 _5089_ (.A(net338),
    .B(net296),
    .X(_2573_));
 sky130_fd_sc_hd__a31o_1 _5090_ (.A1(net434),
    .A2(net1818),
    .A3(net295),
    .B1(_2573_),
    .X(_0287_));
 sky130_fd_sc_hd__and2_1 _5091_ (.A(net336),
    .B(net296),
    .X(_2574_));
 sky130_fd_sc_hd__a31o_1 _5092_ (.A1(net438),
    .A2(net1844),
    .A3(net295),
    .B1(_2574_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_1 _5093_ (.A(net333),
    .B(net296),
    .X(_2575_));
 sky130_fd_sc_hd__a31o_1 _5094_ (.A1(net430),
    .A2(net1809),
    .A3(net295),
    .B1(_2575_),
    .X(_0289_));
 sky130_fd_sc_hd__and2_1 _5095_ (.A(net339),
    .B(net296),
    .X(_2576_));
 sky130_fd_sc_hd__a31o_1 _5096_ (.A1(net433),
    .A2(net1727),
    .A3(net295),
    .B1(_2576_),
    .X(_0290_));
 sky130_fd_sc_hd__and2_1 _5097_ (.A(net340),
    .B(net296),
    .X(_2577_));
 sky130_fd_sc_hd__a31o_1 _5098_ (.A1(net436),
    .A2(net1705),
    .A3(net295),
    .B1(_2577_),
    .X(_0291_));
 sky130_fd_sc_hd__and2_1 _5099_ (.A(net335),
    .B(net296),
    .X(_2578_));
 sky130_fd_sc_hd__a31o_1 _5100_ (.A1(net434),
    .A2(net1611),
    .A3(net295),
    .B1(_2578_),
    .X(_0292_));
 sky130_fd_sc_hd__and2_2 _5101_ (.A(_1287_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_2579_));
 sky130_fd_sc_hd__nand2_2 _5102_ (.A(_1287_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2580_));
 sky130_fd_sc_hd__nor2_2 _5103_ (.A(_2544_),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__or2_1 _5104_ (.A(_2544_),
    .B(_2580_),
    .X(_2582_));
 sky130_fd_sc_hd__nor2_1 _5105_ (.A(net460),
    .B(net293),
    .Y(_2583_));
 sky130_fd_sc_hd__nand2_1 _5106_ (.A(net454),
    .B(_2582_),
    .Y(_2584_));
 sky130_fd_sc_hd__a22o_1 _5107_ (.A1(net298),
    .A2(net293),
    .B1(net237),
    .B2(net1155),
    .X(_0323_));
 sky130_fd_sc_hd__o22a_1 _5108_ (.A1(net299),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net895),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _5109_ (.A1(net353),
    .A2(net293),
    .B1(net237),
    .B2(net1131),
    .X(_0325_));
 sky130_fd_sc_hd__o22a_1 _5110_ (.A1(net355),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net1535),
    .X(_0326_));
 sky130_fd_sc_hd__a22o_1 _5111_ (.A1(net356),
    .A2(net293),
    .B1(net237),
    .B2(net1117),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _5112_ (.A1(net354),
    .A2(net293),
    .B1(net237),
    .B2(net1487),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _5113_ (.A1(net352),
    .A2(net292),
    .B1(net236),
    .B2(net1653),
    .X(_0329_));
 sky130_fd_sc_hd__a22o_1 _5114_ (.A1(net351),
    .A2(net293),
    .B1(net237),
    .B2(net1183),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _5115_ (.A1(net358),
    .A2(net293),
    .B1(net237),
    .B2(net1318),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_1 _5116_ (.A1(net359),
    .A2(net293),
    .B1(net237),
    .B2(net1349),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_1 _5117_ (.A1(net357),
    .A2(net292),
    .B1(net236),
    .B2(net1493),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_1 _5118_ (.A1(net361),
    .A2(net292),
    .B1(net236),
    .B2(net1605),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _5119_ (.A1(_1349_),
    .A2(net293),
    .B1(net237),
    .B2(net1483),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _5120_ (.A1(net360),
    .A2(net292),
    .B1(net236),
    .B2(net1300),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _5121_ (.A1(net350),
    .A2(net293),
    .B1(net237),
    .B2(net1181),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _5122_ (.A1(net349),
    .A2(net293),
    .B1(net237),
    .B2(net1363),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _5123_ (.A1(net345),
    .A2(net292),
    .B1(net236),
    .B2(net1555),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _5124_ (.A1(net344),
    .A2(net293),
    .B1(net237),
    .B2(net1167),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _5125_ (.A1(net341),
    .A2(net293),
    .B1(net237),
    .B2(net1473),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _5126_ (.A1(net343),
    .A2(net292),
    .B1(net236),
    .B2(net1049),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _5127_ (.A1(net342),
    .A2(net292),
    .B1(net236),
    .B2(net1435),
    .X(_0343_));
 sky130_fd_sc_hd__a22o_1 _5128_ (.A1(net346),
    .A2(net292),
    .B1(net236),
    .B2(net1312),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_1 _5129_ (.A1(net348),
    .A2(net293),
    .B1(net237),
    .B2(net1194),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _5130_ (.A1(net347),
    .A2(net292),
    .B1(net236),
    .B2(net1557),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _5131_ (.A1(net334),
    .A2(net293),
    .B1(net237),
    .B2(net1507),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _5132_ (.A1(net337),
    .A2(net292),
    .B1(net236),
    .B2(net1583),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _5133_ (.A1(net338),
    .A2(net292),
    .B1(net236),
    .B2(net1353),
    .X(_0349_));
 sky130_fd_sc_hd__a22o_1 _5134_ (.A1(net336),
    .A2(net292),
    .B1(net236),
    .B2(net1543),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _5135_ (.A1(net333),
    .A2(net292),
    .B1(net236),
    .B2(net1579),
    .X(_0351_));
 sky130_fd_sc_hd__a22o_1 _5136_ (.A1(net339),
    .A2(net292),
    .B1(net236),
    .B2(net1260),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _5137_ (.A1(net340),
    .A2(net292),
    .B1(net236),
    .B2(net1137),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _5138_ (.A1(net335),
    .A2(net292),
    .B1(net236),
    .B2(net1335),
    .X(_0354_));
 sky130_fd_sc_hd__and4_4 _5139_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .B(net453),
    .C(_2507_),
    .D(_2508_),
    .X(_2585_));
 sky130_fd_sc_hd__and2_1 _5140_ (.A(net326),
    .B(net324),
    .X(_2586_));
 sky130_fd_sc_hd__nand2_4 _5141_ (.A(net326),
    .B(net323),
    .Y(_2587_));
 sky130_fd_sc_hd__and2_1 _5142_ (.A(net298),
    .B(_2586_),
    .X(_2588_));
 sky130_fd_sc_hd__a31o_1 _5143_ (.A1(net454),
    .A2(net1926),
    .A3(net290),
    .B1(_2588_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _5144_ (.A(net299),
    .B(_2586_),
    .X(_2589_));
 sky130_fd_sc_hd__a31o_1 _5145_ (.A1(net454),
    .A2(net1964),
    .A3(net290),
    .B1(_2589_),
    .X(_0356_));
 sky130_fd_sc_hd__and3_1 _5146_ (.A(net353),
    .B(net326),
    .C(net323),
    .X(_2590_));
 sky130_fd_sc_hd__a31o_1 _5147_ (.A1(_0069_),
    .A2(net1840),
    .A3(net290),
    .B1(_2590_),
    .X(_0357_));
 sky130_fd_sc_hd__or3_1 _5148_ (.A(net464),
    .B(net2101),
    .C(_2586_),
    .X(_2591_));
 sky130_fd_sc_hd__o21a_1 _5149_ (.A1(net355),
    .A2(net290),
    .B1(_2591_),
    .X(_0358_));
 sky130_fd_sc_hd__and3_1 _5150_ (.A(net356),
    .B(net326),
    .C(net323),
    .X(_2592_));
 sky130_fd_sc_hd__a31o_1 _5151_ (.A1(net455),
    .A2(net1894),
    .A3(net290),
    .B1(_2592_),
    .X(_0359_));
 sky130_fd_sc_hd__and3_1 _5152_ (.A(net354),
    .B(net326),
    .C(net323),
    .X(_2593_));
 sky130_fd_sc_hd__a31o_1 _5153_ (.A1(net455),
    .A2(net1986),
    .A3(net290),
    .B1(_2593_),
    .X(_0360_));
 sky130_fd_sc_hd__and3_1 _5154_ (.A(net352),
    .B(net325),
    .C(net322),
    .X(_2594_));
 sky130_fd_sc_hd__a31o_1 _5155_ (.A1(net439),
    .A2(net1916),
    .A3(net291),
    .B1(_2594_),
    .X(_0361_));
 sky130_fd_sc_hd__and3_1 _5156_ (.A(net351),
    .B(net326),
    .C(net323),
    .X(_2595_));
 sky130_fd_sc_hd__a31o_1 _5157_ (.A1(net446),
    .A2(net1994),
    .A3(net290),
    .B1(_2595_),
    .X(_0362_));
 sky130_fd_sc_hd__and3_1 _5158_ (.A(net358),
    .B(net326),
    .C(net323),
    .X(_2596_));
 sky130_fd_sc_hd__a31o_1 _5159_ (.A1(net446),
    .A2(net1953),
    .A3(net290),
    .B1(_2596_),
    .X(_0363_));
 sky130_fd_sc_hd__and3_1 _5160_ (.A(net359),
    .B(net326),
    .C(net324),
    .X(_2597_));
 sky130_fd_sc_hd__a31o_1 _5161_ (.A1(net456),
    .A2(net1731),
    .A3(net290),
    .B1(_2597_),
    .X(_0364_));
 sky130_fd_sc_hd__and3_1 _5162_ (.A(net357),
    .B(net325),
    .C(net322),
    .X(_2598_));
 sky130_fd_sc_hd__a31o_1 _5163_ (.A1(net446),
    .A2(net1908),
    .A3(net291),
    .B1(_2598_),
    .X(_0365_));
 sky130_fd_sc_hd__and3_1 _5164_ (.A(net361),
    .B(net325),
    .C(net321),
    .X(_2599_));
 sky130_fd_sc_hd__a31o_1 _5165_ (.A1(net433),
    .A2(net1850),
    .A3(net291),
    .B1(_2599_),
    .X(_0366_));
 sky130_fd_sc_hd__nor2_1 _5166_ (.A(_1350_),
    .B(net290),
    .Y(_2600_));
 sky130_fd_sc_hd__a31o_1 _5167_ (.A1(net452),
    .A2(net1967),
    .A3(net290),
    .B1(_2600_),
    .X(_0367_));
 sky130_fd_sc_hd__and3_1 _5168_ (.A(net360),
    .B(net325),
    .C(net322),
    .X(_2601_));
 sky130_fd_sc_hd__a31o_1 _5169_ (.A1(net437),
    .A2(net1974),
    .A3(net291),
    .B1(_2601_),
    .X(_0368_));
 sky130_fd_sc_hd__and3_1 _5170_ (.A(net350),
    .B(net326),
    .C(net323),
    .X(_2602_));
 sky130_fd_sc_hd__a31o_1 _5171_ (.A1(net453),
    .A2(net1932),
    .A3(net290),
    .B1(_2602_),
    .X(_0369_));
 sky130_fd_sc_hd__and3_1 _5172_ (.A(net349),
    .B(net326),
    .C(net323),
    .X(_2603_));
 sky130_fd_sc_hd__a31o_1 _5173_ (.A1(net448),
    .A2(net1822),
    .A3(net290),
    .B1(_2603_),
    .X(_0370_));
 sky130_fd_sc_hd__and3_1 _5174_ (.A(net345),
    .B(net325),
    .C(_2585_),
    .X(_2604_));
 sky130_fd_sc_hd__a31o_1 _5175_ (.A1(net445),
    .A2(net1783),
    .A3(net291),
    .B1(_2604_),
    .X(_0371_));
 sky130_fd_sc_hd__and3_1 _5176_ (.A(net344),
    .B(net326),
    .C(net323),
    .X(_2605_));
 sky130_fd_sc_hd__a31o_1 _5177_ (.A1(net448),
    .A2(net1834),
    .A3(net290),
    .B1(_2605_),
    .X(_0372_));
 sky130_fd_sc_hd__and3_1 _5178_ (.A(net341),
    .B(net326),
    .C(net324),
    .X(_2606_));
 sky130_fd_sc_hd__a31o_1 _5179_ (.A1(net455),
    .A2(net1980),
    .A3(_2587_),
    .B1(_2606_),
    .X(_0373_));
 sky130_fd_sc_hd__and3_1 _5180_ (.A(net343),
    .B(net325),
    .C(net322),
    .X(_2607_));
 sky130_fd_sc_hd__a31o_1 _5181_ (.A1(net437),
    .A2(net1918),
    .A3(net291),
    .B1(_2607_),
    .X(_0374_));
 sky130_fd_sc_hd__and3_1 _5182_ (.A(net342),
    .B(net325),
    .C(net321),
    .X(_2608_));
 sky130_fd_sc_hd__a31o_1 _5183_ (.A1(net436),
    .A2(net1999),
    .A3(net291),
    .B1(_2608_),
    .X(_0375_));
 sky130_fd_sc_hd__and3_1 _5184_ (.A(net346),
    .B(net325),
    .C(net322),
    .X(_2609_));
 sky130_fd_sc_hd__a31o_1 _5185_ (.A1(net437),
    .A2(net1830),
    .A3(net291),
    .B1(_2609_),
    .X(_0376_));
 sky130_fd_sc_hd__and3_1 _5186_ (.A(net348),
    .B(net326),
    .C(net323),
    .X(_2610_));
 sky130_fd_sc_hd__a31o_1 _5187_ (.A1(net445),
    .A2(net1940),
    .A3(net290),
    .B1(_2610_),
    .X(_0377_));
 sky130_fd_sc_hd__and3_1 _5188_ (.A(net347),
    .B(net325),
    .C(net321),
    .X(_2611_));
 sky130_fd_sc_hd__a31o_1 _5189_ (.A1(net434),
    .A2(net1969),
    .A3(net291),
    .B1(_2611_),
    .X(_0378_));
 sky130_fd_sc_hd__and3_1 _5190_ (.A(net334),
    .B(net326),
    .C(net324),
    .X(_2612_));
 sky130_fd_sc_hd__a31o_1 _5191_ (.A1(net456),
    .A2(net1951),
    .A3(net290),
    .B1(_2612_),
    .X(_0379_));
 sky130_fd_sc_hd__and3_1 _5192_ (.A(net337),
    .B(net325),
    .C(net321),
    .X(_2613_));
 sky130_fd_sc_hd__a31o_1 _5193_ (.A1(net433),
    .A2(net1874),
    .A3(net291),
    .B1(_2613_),
    .X(_0380_));
 sky130_fd_sc_hd__and3_1 _5194_ (.A(net338),
    .B(net325),
    .C(net321),
    .X(_2614_));
 sky130_fd_sc_hd__a31o_1 _5195_ (.A1(net434),
    .A2(net1928),
    .A3(net291),
    .B1(_2614_),
    .X(_0381_));
 sky130_fd_sc_hd__and3_1 _5196_ (.A(net336),
    .B(net325),
    .C(net322),
    .X(_2615_));
 sky130_fd_sc_hd__a31o_1 _5197_ (.A1(net439),
    .A2(net1938),
    .A3(net291),
    .B1(_2615_),
    .X(_0382_));
 sky130_fd_sc_hd__and3_1 _5198_ (.A(net333),
    .B(net325),
    .C(net321),
    .X(_2616_));
 sky130_fd_sc_hd__a31o_1 _5199_ (.A1(net433),
    .A2(net1739),
    .A3(net291),
    .B1(_2616_),
    .X(_0383_));
 sky130_fd_sc_hd__and3_1 _5200_ (.A(net339),
    .B(net325),
    .C(net321),
    .X(_2617_));
 sky130_fd_sc_hd__a31o_1 _5201_ (.A1(net433),
    .A2(net1978),
    .A3(net291),
    .B1(_2617_),
    .X(_0384_));
 sky130_fd_sc_hd__and3_1 _5202_ (.A(net340),
    .B(net325),
    .C(net322),
    .X(_2618_));
 sky130_fd_sc_hd__a31o_1 _5203_ (.A1(net436),
    .A2(net1992),
    .A3(net291),
    .B1(_2618_),
    .X(_0385_));
 sky130_fd_sc_hd__and3_1 _5204_ (.A(net335),
    .B(net325),
    .C(net321),
    .X(_2619_));
 sky130_fd_sc_hd__a31o_1 _5205_ (.A1(net433),
    .A2(net1860),
    .A3(net291),
    .B1(_2619_),
    .X(_0386_));
 sky130_fd_sc_hd__and4_2 _5206_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .D(net454),
    .X(_2620_));
 sky130_fd_sc_hd__and2_2 _5207_ (.A(net326),
    .B(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__nand2_1 _5208_ (.A(net326),
    .B(_2620_),
    .Y(_2622_));
 sky130_fd_sc_hd__nor2_2 _5209_ (.A(net464),
    .B(net289),
    .Y(_2623_));
 sky130_fd_sc_hd__nand2_1 _5210_ (.A(net454),
    .B(_2622_),
    .Y(_2624_));
 sky130_fd_sc_hd__o22a_1 _5211_ (.A1(net298),
    .A2(_2622_),
    .B1(_2624_),
    .B2(net877),
    .X(_0387_));
 sky130_fd_sc_hd__o22a_1 _5212_ (.A1(net299),
    .A2(_2622_),
    .B1(_2624_),
    .B2(net881),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _5213_ (.A1(net353),
    .A2(net289),
    .B1(net235),
    .B2(net1051),
    .X(_0389_));
 sky130_fd_sc_hd__o22a_1 _5214_ (.A1(net355),
    .A2(_2622_),
    .B1(_2624_),
    .B2(net1133),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _5215_ (.A1(net356),
    .A2(net289),
    .B1(net235),
    .B2(net1680),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _5216_ (.A1(net354),
    .A2(net289),
    .B1(net235),
    .B2(net1240),
    .X(_0392_));
 sky130_fd_sc_hd__a22o_1 _5217_ (.A1(net352),
    .A2(net288),
    .B1(net234),
    .B2(net1467),
    .X(_0393_));
 sky130_fd_sc_hd__a22o_1 _5218_ (.A1(net351),
    .A2(net289),
    .B1(net235),
    .B2(net1643),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_1 _5219_ (.A1(net358),
    .A2(net289),
    .B1(net235),
    .B2(net1270),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _5220_ (.A1(net359),
    .A2(net289),
    .B1(net235),
    .B2(net1163),
    .X(_0396_));
 sky130_fd_sc_hd__a22o_1 _5221_ (.A1(net357),
    .A2(net288),
    .B1(net234),
    .B2(net1222),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _5222_ (.A1(net361),
    .A2(net288),
    .B1(net234),
    .B2(net1383),
    .X(_0398_));
 sky130_fd_sc_hd__a22o_1 _5223_ (.A1(_1349_),
    .A2(net289),
    .B1(net235),
    .B2(net1304),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_1 _5224_ (.A1(net360),
    .A2(net288),
    .B1(net234),
    .B2(net1125),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_1 _5225_ (.A1(net350),
    .A2(net289),
    .B1(net235),
    .B2(net1218),
    .X(_0401_));
 sky130_fd_sc_hd__a22o_1 _5226_ (.A1(net349),
    .A2(net289),
    .B1(net235),
    .B2(net1087),
    .X(_0402_));
 sky130_fd_sc_hd__a22o_1 _5227_ (.A1(net345),
    .A2(net288),
    .B1(net234),
    .B2(net1664),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _5228_ (.A1(net344),
    .A2(net289),
    .B1(net235),
    .B2(net1505),
    .X(_0404_));
 sky130_fd_sc_hd__a22o_1 _5229_ (.A1(net341),
    .A2(net289),
    .B1(net235),
    .B2(net1258),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _5230_ (.A1(net343),
    .A2(net288),
    .B1(net234),
    .B2(net1113),
    .X(_0406_));
 sky130_fd_sc_hd__a22o_1 _5231_ (.A1(net342),
    .A2(net288),
    .B1(net234),
    .B2(net1674),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _5232_ (.A1(net346),
    .A2(net288),
    .B1(net234),
    .B2(net1684),
    .X(_0408_));
 sky130_fd_sc_hd__a22o_1 _5233_ (.A1(net348),
    .A2(net289),
    .B1(net235),
    .B2(net1595),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _5234_ (.A1(net347),
    .A2(net288),
    .B1(net234),
    .B2(net1629),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_1 _5235_ (.A1(net334),
    .A2(net289),
    .B1(net235),
    .B2(net1387),
    .X(_0411_));
 sky130_fd_sc_hd__a22o_1 _5236_ (.A1(net337),
    .A2(net288),
    .B1(net234),
    .B2(net1858),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _5237_ (.A1(net338),
    .A2(net288),
    .B1(net234),
    .B2(net1165),
    .X(_0413_));
 sky130_fd_sc_hd__a22o_1 _5238_ (.A1(net336),
    .A2(net288),
    .B1(net234),
    .B2(net1371),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _5239_ (.A1(net333),
    .A2(net288),
    .B1(net234),
    .B2(net1577),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _5240_ (.A1(net339),
    .A2(net288),
    .B1(net234),
    .B2(net1499),
    .X(_0416_));
 sky130_fd_sc_hd__a22o_1 _5241_ (.A1(net340),
    .A2(net288),
    .B1(net234),
    .B2(net1041),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _5242_ (.A1(net335),
    .A2(net288),
    .B1(net234),
    .B2(net1039),
    .X(_0418_));
 sky130_fd_sc_hd__nor2_2 _5243_ (.A(_1287_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2625_));
 sky130_fd_sc_hd__or2_1 _5244_ (.A(_1287_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_2626_));
 sky130_fd_sc_hd__and2_1 _5245_ (.A(net323),
    .B(net320),
    .X(_2627_));
 sky130_fd_sc_hd__nand2_4 _5246_ (.A(net323),
    .B(net320),
    .Y(_2628_));
 sky130_fd_sc_hd__and2_1 _5247_ (.A(net298),
    .B(_2627_),
    .X(_2629_));
 sky130_fd_sc_hd__a31o_1 _5248_ (.A1(net447),
    .A2(net1984),
    .A3(net287),
    .B1(_2629_),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _5249_ (.A(net299),
    .B(_2627_),
    .X(_2630_));
 sky130_fd_sc_hd__a31o_1 _5250_ (.A1(net447),
    .A2(net1976),
    .A3(net287),
    .B1(_2630_),
    .X(_0420_));
 sky130_fd_sc_hd__or3_1 _5251_ (.A(net464),
    .B(net2111),
    .C(_2627_),
    .X(_2631_));
 sky130_fd_sc_hd__o21a_1 _5252_ (.A1(net353),
    .A2(net287),
    .B1(_2631_),
    .X(_0421_));
 sky130_fd_sc_hd__and3_1 _5253_ (.A(net355),
    .B(net324),
    .C(net320),
    .X(_2632_));
 sky130_fd_sc_hd__a31o_1 _5254_ (.A1(net456),
    .A2(net1944),
    .A3(net287),
    .B1(_2632_),
    .X(_0422_));
 sky130_fd_sc_hd__and3_1 _5255_ (.A(net356),
    .B(net324),
    .C(net320),
    .X(_2633_));
 sky130_fd_sc_hd__a31o_1 _5256_ (.A1(net455),
    .A2(net1982),
    .A3(net287),
    .B1(_2633_),
    .X(_0423_));
 sky130_fd_sc_hd__and3_1 _5257_ (.A(net354),
    .B(net324),
    .C(net320),
    .X(_2634_));
 sky130_fd_sc_hd__a31o_1 _5258_ (.A1(net452),
    .A2(net1775),
    .A3(net287),
    .B1(_2634_),
    .X(_0424_));
 sky130_fd_sc_hd__and3_1 _5259_ (.A(net352),
    .B(net322),
    .C(net319),
    .X(_2635_));
 sky130_fd_sc_hd__a31o_1 _5260_ (.A1(net439),
    .A2(net1692),
    .A3(net287),
    .B1(_2635_),
    .X(_0425_));
 sky130_fd_sc_hd__and3_1 _5261_ (.A(net351),
    .B(_2585_),
    .C(net319),
    .X(_2636_));
 sky130_fd_sc_hd__a31o_1 _5262_ (.A1(net445),
    .A2(net1888),
    .A3(net286),
    .B1(_2636_),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _5263_ (.A(net358),
    .B(net322),
    .C(net319),
    .X(_2637_));
 sky130_fd_sc_hd__a31o_1 _5264_ (.A1(net446),
    .A2(net1971),
    .A3(net286),
    .B1(_2637_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _5265_ (.A(net359),
    .B(net324),
    .C(net320),
    .X(_2638_));
 sky130_fd_sc_hd__a31o_1 _5266_ (.A1(net455),
    .A2(net1666),
    .A3(net287),
    .B1(_2638_),
    .X(_0428_));
 sky130_fd_sc_hd__and3_1 _5267_ (.A(net357),
    .B(net322),
    .C(net319),
    .X(_2639_));
 sky130_fd_sc_hd__a31o_1 _5268_ (.A1(net445),
    .A2(net1936),
    .A3(net286),
    .B1(_2639_),
    .X(_0429_));
 sky130_fd_sc_hd__and3_1 _5269_ (.A(net361),
    .B(net321),
    .C(net319),
    .X(_2640_));
 sky130_fd_sc_hd__a31o_1 _5270_ (.A1(net441),
    .A2(net1962),
    .A3(net286),
    .B1(_2640_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_1 _5271_ (.A(_1350_),
    .B(net287),
    .Y(_2641_));
 sky130_fd_sc_hd__a31o_1 _5272_ (.A1(net452),
    .A2(net1862),
    .A3(net287),
    .B1(_2641_),
    .X(_0431_));
 sky130_fd_sc_hd__and3_1 _5273_ (.A(net360),
    .B(net322),
    .C(net319),
    .X(_2642_));
 sky130_fd_sc_hd__a31o_1 _5274_ (.A1(net437),
    .A2(net1898),
    .A3(net287),
    .B1(_2642_),
    .X(_0432_));
 sky130_fd_sc_hd__and3_1 _5275_ (.A(net350),
    .B(net323),
    .C(net320),
    .X(_2643_));
 sky130_fd_sc_hd__a31o_1 _5276_ (.A1(net451),
    .A2(net1761),
    .A3(net287),
    .B1(_2643_),
    .X(_0433_));
 sky130_fd_sc_hd__and3_1 _5277_ (.A(net349),
    .B(net324),
    .C(net320),
    .X(_2644_));
 sky130_fd_sc_hd__a31o_1 _5278_ (.A1(net451),
    .A2(net1892),
    .A3(net287),
    .B1(_2644_),
    .X(_0434_));
 sky130_fd_sc_hd__and3_1 _5279_ (.A(net345),
    .B(_2585_),
    .C(net320),
    .X(_2645_));
 sky130_fd_sc_hd__a31o_1 _5280_ (.A1(net445),
    .A2(net1878),
    .A3(net286),
    .B1(_2645_),
    .X(_0435_));
 sky130_fd_sc_hd__and3_1 _5281_ (.A(net344),
    .B(net323),
    .C(net320),
    .X(_2646_));
 sky130_fd_sc_hd__a31o_1 _5282_ (.A1(net453),
    .A2(net1884),
    .A3(net287),
    .B1(_2646_),
    .X(_0436_));
 sky130_fd_sc_hd__and3_1 _5283_ (.A(net341),
    .B(net324),
    .C(_2625_),
    .X(_2647_));
 sky130_fd_sc_hd__a31o_1 _5284_ (.A1(net455),
    .A2(net1824),
    .A3(_2628_),
    .B1(_2647_),
    .X(_0437_));
 sky130_fd_sc_hd__and3_1 _5285_ (.A(net343),
    .B(net322),
    .C(net319),
    .X(_2648_));
 sky130_fd_sc_hd__a31o_1 _5286_ (.A1(net438),
    .A2(net1910),
    .A3(net286),
    .B1(_2648_),
    .X(_0438_));
 sky130_fd_sc_hd__and3_1 _5287_ (.A(net342),
    .B(net322),
    .C(net319),
    .X(_2649_));
 sky130_fd_sc_hd__a31o_1 _5288_ (.A1(net436),
    .A2(net1789),
    .A3(net286),
    .B1(_2649_),
    .X(_0439_));
 sky130_fd_sc_hd__and3_1 _5289_ (.A(net346),
    .B(net321),
    .C(net319),
    .X(_2650_));
 sky130_fd_sc_hd__a31o_1 _5290_ (.A1(net436),
    .A2(net1996),
    .A3(net286),
    .B1(_2650_),
    .X(_0440_));
 sky130_fd_sc_hd__and3_1 _5291_ (.A(net348),
    .B(net323),
    .C(net320),
    .X(_2651_));
 sky130_fd_sc_hd__a31o_1 _5292_ (.A1(net447),
    .A2(net1852),
    .A3(net287),
    .B1(_2651_),
    .X(_0441_));
 sky130_fd_sc_hd__and3_1 _5293_ (.A(net347),
    .B(net321),
    .C(net319),
    .X(_2652_));
 sky130_fd_sc_hd__a31o_1 _5294_ (.A1(net434),
    .A2(net1922),
    .A3(net286),
    .B1(_2652_),
    .X(_0442_));
 sky130_fd_sc_hd__and3_1 _5295_ (.A(net334),
    .B(net324),
    .C(net320),
    .X(_2653_));
 sky130_fd_sc_hd__a31o_1 _5296_ (.A1(net455),
    .A2(net1791),
    .A3(_2628_),
    .B1(_2653_),
    .X(_0443_));
 sky130_fd_sc_hd__and3_1 _5297_ (.A(net337),
    .B(net321),
    .C(net319),
    .X(_2654_));
 sky130_fd_sc_hd__a31o_1 _5298_ (.A1(net433),
    .A2(net1930),
    .A3(net286),
    .B1(_2654_),
    .X(_0444_));
 sky130_fd_sc_hd__and3_1 _5299_ (.A(net338),
    .B(net321),
    .C(net319),
    .X(_2655_));
 sky130_fd_sc_hd__a31o_1 _5300_ (.A1(net434),
    .A2(net1856),
    .A3(net286),
    .B1(_2655_),
    .X(_0445_));
 sky130_fd_sc_hd__and3_1 _5301_ (.A(net336),
    .B(net322),
    .C(net320),
    .X(_2656_));
 sky130_fd_sc_hd__a31o_1 _5302_ (.A1(net445),
    .A2(net1799),
    .A3(net286),
    .B1(_2656_),
    .X(_0446_));
 sky130_fd_sc_hd__and3_1 _5303_ (.A(net333),
    .B(net321),
    .C(net319),
    .X(_2657_));
 sky130_fd_sc_hd__a31o_1 _5304_ (.A1(net441),
    .A2(net1771),
    .A3(net286),
    .B1(_2657_),
    .X(_0447_));
 sky130_fd_sc_hd__and3_1 _5305_ (.A(net339),
    .B(net321),
    .C(net319),
    .X(_2658_));
 sky130_fd_sc_hd__a31o_1 _5306_ (.A1(net433),
    .A2(net1900),
    .A3(net286),
    .B1(_2658_),
    .X(_0448_));
 sky130_fd_sc_hd__and3_1 _5307_ (.A(net340),
    .B(net322),
    .C(net319),
    .X(_2659_));
 sky130_fd_sc_hd__a31o_1 _5308_ (.A1(net436),
    .A2(net1960),
    .A3(net286),
    .B1(_2659_),
    .X(_0449_));
 sky130_fd_sc_hd__and3_1 _5309_ (.A(net335),
    .B(net321),
    .C(net319),
    .X(_2660_));
 sky130_fd_sc_hd__a31o_1 _5310_ (.A1(net437),
    .A2(net1957),
    .A3(net286),
    .B1(_2660_),
    .X(_0450_));
 sky130_fd_sc_hd__and2b_2 _5311_ (.A_N(_2507_),
    .B(_2620_),
    .X(_2661_));
 sky130_fd_sc_hd__nand2b_1 _5312_ (.A_N(_2507_),
    .B(_2620_),
    .Y(_2662_));
 sky130_fd_sc_hd__nor2_2 _5313_ (.A(net460),
    .B(net318),
    .Y(_2663_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(net454),
    .B(_2662_),
    .Y(_2664_));
 sky130_fd_sc_hd__o22a_1 _5315_ (.A1(net298),
    .A2(_2662_),
    .B1(_2664_),
    .B2(net970),
    .X(_0451_));
 sky130_fd_sc_hd__o22a_1 _5316_ (.A1(net299),
    .A2(_2662_),
    .B1(_2664_),
    .B2(net1719),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _5317_ (.A1(net353),
    .A2(net318),
    .B1(net285),
    .B2(net1682),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _5318_ (.A1(net355),
    .A2(net318),
    .B1(net285),
    .B2(net1057),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _5319_ (.A1(net356),
    .A2(net318),
    .B1(net285),
    .B2(net1306),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _5320_ (.A1(net354),
    .A2(net318),
    .B1(net285),
    .B2(net1149),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _5321_ (.A1(net352),
    .A2(net317),
    .B1(net284),
    .B2(net983),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _5322_ (.A1(net351),
    .A2(net318),
    .B1(net285),
    .B2(net1575),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(net358),
    .A2(net317),
    .B1(net284),
    .B2(net1459),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _5324_ (.A1(net359),
    .A2(net318),
    .B1(net285),
    .B2(net1028),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _5325_ (.A1(net357),
    .A2(net317),
    .B1(net284),
    .B2(net1461),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _5326_ (.A1(net361),
    .A2(net317),
    .B1(net284),
    .B2(net1037),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _5327_ (.A1(_1349_),
    .A2(net318),
    .B1(net285),
    .B2(net1471),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _5328_ (.A1(net360),
    .A2(net317),
    .B1(net284),
    .B2(net1397),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _5329_ (.A1(net350),
    .A2(net318),
    .B1(net285),
    .B2(net1097),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _5330_ (.A1(net349),
    .A2(net318),
    .B1(net285),
    .B2(net1014),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(net345),
    .A2(net318),
    .B1(net285),
    .B2(net1296),
    .X(_0467_));
 sky130_fd_sc_hd__a22o_1 _5332_ (.A1(net344),
    .A2(net318),
    .B1(net285),
    .B2(net1161),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _5333_ (.A1(net341),
    .A2(net318),
    .B1(net285),
    .B2(net1121),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _5334_ (.A1(net343),
    .A2(net317),
    .B1(net284),
    .B2(net1331),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _5335_ (.A1(net342),
    .A2(net317),
    .B1(net284),
    .B2(net1071),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _5336_ (.A1(net346),
    .A2(net317),
    .B1(net284),
    .B2(net1298),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _5337_ (.A1(net348),
    .A2(net318),
    .B1(net285),
    .B2(net1395),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _5338_ (.A1(net347),
    .A2(net317),
    .B1(net284),
    .B2(net1216),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _5339_ (.A1(net334),
    .A2(net318),
    .B1(net285),
    .B2(net1145),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _5340_ (.A1(net337),
    .A2(net317),
    .B1(net284),
    .B2(net1405),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _5341_ (.A1(net338),
    .A2(net317),
    .B1(net284),
    .B2(net1729),
    .X(_0477_));
 sky130_fd_sc_hd__a22o_1 _5342_ (.A1(net336),
    .A2(net317),
    .B1(net284),
    .B2(net1355),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _5343_ (.A1(net333),
    .A2(net317),
    .B1(net284),
    .B2(net1246),
    .X(_0479_));
 sky130_fd_sc_hd__a22o_1 _5344_ (.A1(net339),
    .A2(net317),
    .B1(net284),
    .B2(net961),
    .X(_0480_));
 sky130_fd_sc_hd__a22o_1 _5345_ (.A1(net340),
    .A2(net317),
    .B1(net284),
    .B2(net985),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _5346_ (.A1(net335),
    .A2(net317),
    .B1(net284),
    .B2(net1288),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _5347_ (.A(_0067_),
    .B(_2474_),
    .Y(_2665_));
 sky130_fd_sc_hd__a21o_1 _5348_ (.A1(_1278_),
    .A2(net2148),
    .B1(_2477_),
    .X(_2666_));
 sky130_fd_sc_hd__a32o_1 _5349_ (.A1(net2119),
    .A2(net2148),
    .A3(_2464_),
    .B1(_2665_),
    .B2(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__a21boi_1 _5350_ (.A1(_2470_),
    .A2(_2667_),
    .B1_N(_2497_),
    .Y(_2668_));
 sky130_fd_sc_hd__o211a_1 _5351_ (.A1(_2487_),
    .A2(_2668_),
    .B1(_2491_),
    .C1(net176),
    .X(_0483_));
 sky130_fd_sc_hd__and2_2 _5352_ (.A(net426),
    .B(net179),
    .X(_0484_));
 sky130_fd_sc_hd__nor2_2 _5353_ (.A(_1279_),
    .B(net162),
    .Y(_0485_));
 sky130_fd_sc_hd__nor2_1 _5354_ (.A(_1278_),
    .B(net162),
    .Y(_0486_));
 sky130_fd_sc_hd__and2_1 _5355_ (.A(net2129),
    .B(net447),
    .X(_0487_));
 sky130_fd_sc_hd__and2_1 _5356_ (.A(net2086),
    .B(net447),
    .X(_0488_));
 sky130_fd_sc_hd__and2_1 _5357_ (.A(net2220),
    .B(net448),
    .X(_0489_));
 sky130_fd_sc_hd__and2_1 _5358_ (.A(net1701),
    .B(net451),
    .X(_0490_));
 sky130_fd_sc_hd__and2_1 _5359_ (.A(net1007),
    .B(net450),
    .X(_0491_));
 sky130_fd_sc_hd__and2_1 _5360_ (.A(net2100),
    .B(net451),
    .X(_0492_));
 sky130_fd_sc_hd__and2_1 _5361_ (.A(net2146),
    .B(net446),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _5362_ (.A(net2210),
    .B(net443),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _5363_ (.A(net2192),
    .B(net444),
    .X(_0495_));
 sky130_fd_sc_hd__and2_1 _5364_ (.A(net860),
    .B(net451),
    .X(_0496_));
 sky130_fd_sc_hd__and2_1 _5365_ (.A(net2087),
    .B(net435),
    .X(_0497_));
 sky130_fd_sc_hd__and2_1 _5366_ (.A(net2166),
    .B(net429),
    .X(_0498_));
 sky130_fd_sc_hd__and2_1 _5367_ (.A(net1655),
    .B(net450),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _5368_ (.A(net2187),
    .B(net438),
    .X(_0500_));
 sky130_fd_sc_hd__and2_1 _5369_ (.A(net2133),
    .B(net451),
    .X(_0501_));
 sky130_fd_sc_hd__and2_1 _5370_ (.A(net2092),
    .B(net442),
    .X(_0502_));
 sky130_fd_sc_hd__and2_1 _5371_ (.A(net2223),
    .B(net446),
    .X(_0503_));
 sky130_fd_sc_hd__and2_1 _5372_ (.A(net2149),
    .B(net448),
    .X(_0504_));
 sky130_fd_sc_hd__and2_1 _5373_ (.A(net2012),
    .B(net453),
    .X(_0505_));
 sky130_fd_sc_hd__and2_1 _5374_ (.A(net2198),
    .B(net438),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _5375_ (.A(net2023),
    .B(net433),
    .X(_0507_));
 sky130_fd_sc_hd__and2_1 _5376_ (.A(net2032),
    .B(net431),
    .X(_0508_));
 sky130_fd_sc_hd__and2_1 _5377_ (.A(net2058),
    .B(net432),
    .X(_0509_));
 sky130_fd_sc_hd__and2_1 _5378_ (.A(net969),
    .B(net432),
    .X(_0510_));
 sky130_fd_sc_hd__and2_1 _5379_ (.A(net2103),
    .B(net436),
    .X(_0511_));
 sky130_fd_sc_hd__and2_1 _5380_ (.A(net537),
    .B(net432),
    .X(_0512_));
 sky130_fd_sc_hd__and2_1 _5381_ (.A(net2024),
    .B(net431),
    .X(_0513_));
 sky130_fd_sc_hd__and2_1 _5382_ (.A(net2143),
    .B(net437),
    .X(_0514_));
 sky130_fd_sc_hd__and2_1 _5383_ (.A(net1704),
    .B(net430),
    .X(_0515_));
 sky130_fd_sc_hd__and2_1 _5384_ (.A(net2186),
    .B(net430),
    .X(_0516_));
 sky130_fd_sc_hd__and2_1 _5385_ (.A(net2125),
    .B(net435),
    .X(_0517_));
 sky130_fd_sc_hd__and2_1 _5386_ (.A(net2163),
    .B(net431),
    .X(_0518_));
 sky130_fd_sc_hd__and2_1 _5387_ (.A(net447),
    .B(net1541),
    .X(_0519_));
 sky130_fd_sc_hd__and2_1 _5388_ (.A(net447),
    .B(net808),
    .X(_0520_));
 sky130_fd_sc_hd__and2_1 _5389_ (.A(net453),
    .B(net784),
    .X(_0521_));
 sky130_fd_sc_hd__and2_1 _5390_ (.A(net451),
    .B(net590),
    .X(_0522_));
 sky130_fd_sc_hd__and2_1 _5391_ (.A(net450),
    .B(net704),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _5392_ (.A(net449),
    .B(net660),
    .X(_0524_));
 sky130_fd_sc_hd__and2_1 _5393_ (.A(net448),
    .B(net640),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _5394_ (.A(net443),
    .B(net632),
    .X(_0526_));
 sky130_fd_sc_hd__and2_1 _5395_ (.A(net442),
    .B(net744),
    .X(_0527_));
 sky130_fd_sc_hd__and2_1 _5396_ (.A(net450),
    .B(net780),
    .X(_0528_));
 sky130_fd_sc_hd__and2_1 _5397_ (.A(net435),
    .B(net592),
    .X(_0529_));
 sky130_fd_sc_hd__and2_1 _5398_ (.A(net429),
    .B(net720),
    .X(_0530_));
 sky130_fd_sc_hd__and2_1 _5399_ (.A(net449),
    .B(net738),
    .X(_0531_));
 sky130_fd_sc_hd__and2_1 _5400_ (.A(net443),
    .B(net600),
    .X(_0532_));
 sky130_fd_sc_hd__and2_1 _5401_ (.A(net449),
    .B(net724),
    .X(_0533_));
 sky130_fd_sc_hd__and2_1 _5402_ (.A(net442),
    .B(net762),
    .X(_0534_));
 sky130_fd_sc_hd__and2_1 _5403_ (.A(net444),
    .B(net553),
    .X(_0535_));
 sky130_fd_sc_hd__and2_1 _5404_ (.A(net448),
    .B(net648),
    .X(_0536_));
 sky130_fd_sc_hd__and2_1 _5405_ (.A(net453),
    .B(net680),
    .X(_0537_));
 sky130_fd_sc_hd__and2_1 _5406_ (.A(net438),
    .B(net690),
    .X(_0538_));
 sky130_fd_sc_hd__and2_1 _5407_ (.A(net432),
    .B(net619),
    .X(_0539_));
 sky130_fd_sc_hd__and2_1 _5408_ (.A(net431),
    .B(net602),
    .X(_0540_));
 sky130_fd_sc_hd__and2_1 _5409_ (.A(net430),
    .B(net789),
    .X(_0541_));
 sky130_fd_sc_hd__and2_1 _5410_ (.A(net432),
    .B(net662),
    .X(_0542_));
 sky130_fd_sc_hd__and2_1 _5411_ (.A(net432),
    .B(net636),
    .X(_0543_));
 sky130_fd_sc_hd__and2_1 _5412_ (.A(net432),
    .B(net654),
    .X(_0544_));
 sky130_fd_sc_hd__and2_1 _5413_ (.A(net431),
    .B(net569),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _5414_ (.A(net431),
    .B(net957),
    .X(_0546_));
 sky130_fd_sc_hd__and2_1 _5415_ (.A(net430),
    .B(net638),
    .X(_0547_));
 sky130_fd_sc_hd__and2_1 _5416_ (.A(net429),
    .B(net598),
    .X(_0548_));
 sky130_fd_sc_hd__and2_1 _5417_ (.A(net429),
    .B(net748),
    .X(_0549_));
 sky130_fd_sc_hd__and2_1 _5418_ (.A(net431),
    .B(net714),
    .X(_0550_));
 sky130_fd_sc_hd__and2_1 _5419_ (.A(net453),
    .B(net623),
    .X(_0551_));
 sky130_fd_sc_hd__and2_1 _5420_ (.A(net451),
    .B(net573),
    .X(_0552_));
 sky130_fd_sc_hd__and2_1 _5421_ (.A(net450),
    .B(net760),
    .X(_0553_));
 sky130_fd_sc_hd__and2_1 _5422_ (.A(net449),
    .B(net686),
    .X(_0554_));
 sky130_fd_sc_hd__and2_1 _5423_ (.A(net448),
    .B(net664),
    .X(_0555_));
 sky130_fd_sc_hd__and2_1 _5424_ (.A(net442),
    .B(net625),
    .X(_0556_));
 sky130_fd_sc_hd__and2_1 _5425_ (.A(net442),
    .B(net615),
    .X(_0557_));
 sky130_fd_sc_hd__and2_1 _5426_ (.A(net449),
    .B(net764),
    .X(_0558_));
 sky130_fd_sc_hd__and2_1 _5427_ (.A(net435),
    .B(net583),
    .X(_0559_));
 sky130_fd_sc_hd__and2_1 _5428_ (.A(net429),
    .B(net688),
    .X(_0560_));
 sky130_fd_sc_hd__and2_1 _5429_ (.A(net450),
    .B(net670),
    .X(_0561_));
 sky130_fd_sc_hd__and2_1 _5430_ (.A(net446),
    .B(net728),
    .X(_0562_));
 sky130_fd_sc_hd__and2_1 _5431_ (.A(net449),
    .B(net652),
    .X(_0563_));
 sky130_fd_sc_hd__and2_1 _5432_ (.A(net442),
    .B(net740),
    .X(_0564_));
 sky130_fd_sc_hd__and2_1 _5433_ (.A(net443),
    .B(net547),
    .X(_0565_));
 sky130_fd_sc_hd__and2_1 _5434_ (.A(net448),
    .B(net678),
    .X(_0566_));
 sky130_fd_sc_hd__and2_1 _5435_ (.A(net453),
    .B(net716),
    .X(_0567_));
 sky130_fd_sc_hd__and2_1 _5436_ (.A(net438),
    .B(net746),
    .X(_0568_));
 sky130_fd_sc_hd__and2_1 _5437_ (.A(net432),
    .B(net712),
    .X(_0569_));
 sky130_fd_sc_hd__and2_1 _5438_ (.A(net431),
    .B(net710),
    .X(_0570_));
 sky130_fd_sc_hd__and2_1 _5439_ (.A(net430),
    .B(net545),
    .X(_0571_));
 sky130_fd_sc_hd__and2_1 _5440_ (.A(net432),
    .B(net702),
    .X(_0572_));
 sky130_fd_sc_hd__and2_1 _5441_ (.A(net436),
    .B(net734),
    .X(_0573_));
 sky130_fd_sc_hd__and2_1 _5442_ (.A(net432),
    .B(net672),
    .X(_0574_));
 sky130_fd_sc_hd__and2_1 _5443_ (.A(net431),
    .B(net750),
    .X(_0575_));
 sky130_fd_sc_hd__and2_1 _5444_ (.A(net441),
    .B(net1513),
    .X(_0576_));
 sky130_fd_sc_hd__and2_1 _5445_ (.A(net430),
    .B(net621),
    .X(_0577_));
 sky130_fd_sc_hd__and2_1 _5446_ (.A(net429),
    .B(net730),
    .X(_0578_));
 sky130_fd_sc_hd__and2_1 _5447_ (.A(net429),
    .B(net766),
    .X(_0579_));
 sky130_fd_sc_hd__and2_1 _5448_ (.A(net431),
    .B(net736),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A1(net2104),
    .S(net464),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _5450_ (.A0(net1177),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .S(net464),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _5451_ (.A0(net2117),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .S(net464),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(net2144),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .S(net464),
    .X(_0584_));
 sky130_fd_sc_hd__and2_1 _5453_ (.A(net851),
    .B(net453),
    .X(_0585_));
 sky130_fd_sc_hd__and2_1 _5454_ (.A(net452),
    .B(net698),
    .X(_0586_));
 sky130_fd_sc_hd__and2_1 _5455_ (.A(net452),
    .B(net555),
    .X(_0587_));
 sky130_fd_sc_hd__and2_1 _5456_ (.A(net435),
    .B(net676),
    .X(_0588_));
 sky130_fd_sc_hd__and2_1 _5457_ (.A(net444),
    .B(net2262),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _5458_ (.A(net460),
    .B(_1474_),
    .Y(_0590_));
 sky130_fd_sc_hd__o31a_4 _5459_ (.A1(_1444_),
    .A2(_1445_),
    .A3(_1446_),
    .B1(net446),
    .X(_0591_));
 sky130_fd_sc_hd__nor2_4 _5460_ (.A(net460),
    .B(_1464_),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2_1 _5461_ (.A(net463),
    .B(_1432_),
    .Y(_0593_));
 sky130_fd_sc_hd__nor2_1 _5462_ (.A(net463),
    .B(_1422_),
    .Y(_0594_));
 sky130_fd_sc_hd__nor2_1 _5463_ (.A(net463),
    .B(_1455_),
    .Y(_0595_));
 sky130_fd_sc_hd__and2_1 _5464_ (.A(net442),
    .B(_1485_),
    .X(_0596_));
 sky130_fd_sc_hd__and2_1 _5465_ (.A(net446),
    .B(net2232),
    .X(_0597_));
 sky130_fd_sc_hd__and2_1 _5466_ (.A(net429),
    .B(_1404_),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _5467_ (.A(net461),
    .B(net2085),
    .Y(_0599_));
 sky130_fd_sc_hd__and2_1 _5468_ (.A(net445),
    .B(_1414_),
    .X(_0600_));
 sky130_fd_sc_hd__nor2_1 _5469_ (.A(net457),
    .B(_1376_),
    .Y(_0601_));
 sky130_fd_sc_hd__and2_1 _5470_ (.A(net442),
    .B(_1353_),
    .X(_0602_));
 sky130_fd_sc_hd__and2_2 _5471_ (.A(net439),
    .B(_1386_),
    .X(_0603_));
 sky130_fd_sc_hd__and2_1 _5472_ (.A(net435),
    .B(_1503_),
    .X(_0604_));
 sky130_fd_sc_hd__and2_1 _5473_ (.A(net444),
    .B(_1510_),
    .X(_0605_));
 sky130_fd_sc_hd__nor2_1 _5474_ (.A(net461),
    .B(_1547_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_1 _5475_ (.A(net460),
    .B(_1556_),
    .Y(_0607_));
 sky130_fd_sc_hd__and2_1 _5476_ (.A(net452),
    .B(_1581_),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_1 _5477_ (.A(net460),
    .B(_1563_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _5478_ (.A(net457),
    .B(_1571_),
    .Y(_0610_));
 sky130_fd_sc_hd__nor2_1 _5479_ (.A(net457),
    .B(_1537_),
    .Y(_0611_));
 sky130_fd_sc_hd__and2_1 _5480_ (.A(net452),
    .B(_1521_),
    .X(_0612_));
 sky130_fd_sc_hd__nor2_1 _5481_ (.A(net458),
    .B(_1528_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_1 _5482_ (.A(net464),
    .B(_1644_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _5483_ (.A(net63),
    .B(net550),
    .Y(_0615_));
 sky130_fd_sc_hd__and2_1 _5484_ (.A(net429),
    .B(_1607_),
    .X(_0616_));
 sky130_fd_sc_hd__and2_1 _5485_ (.A(net447),
    .B(_1624_),
    .X(_0617_));
 sky130_fd_sc_hd__and2_1 _5486_ (.A(net429),
    .B(_1653_),
    .X(_0618_));
 sky130_fd_sc_hd__nor2_1 _5487_ (.A(net457),
    .B(net2182),
    .Y(_0619_));
 sky130_fd_sc_hd__and2_1 _5488_ (.A(net447),
    .B(_1590_),
    .X(_0620_));
 sky130_fd_sc_hd__and2_1 _5489_ (.A(net431),
    .B(_1634_),
    .X(_0621_));
 sky130_fd_sc_hd__and2_1 _5490_ (.A(net449),
    .B(net722),
    .X(_0622_));
 sky130_fd_sc_hd__and2_1 _5491_ (.A(net1619),
    .B(net449),
    .X(_0623_));
 sky130_fd_sc_hd__and2_1 _5492_ (.A(net1282),
    .B(net449),
    .X(_0624_));
 sky130_fd_sc_hd__nand3b_2 _5493_ (.A_N(net2254),
    .B(_1693_),
    .C(_1661_),
    .Y(_2669_));
 sky130_fd_sc_hd__or3b_4 _5494_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(net2208),
    .C_N(net2252),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_4 _5495_ (.A(_1698_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__or2_4 _5496_ (.A(_1698_),
    .B(_2670_),
    .X(_2672_));
 sky130_fd_sc_hd__nor2_4 _5497_ (.A(_1700_),
    .B(_1703_),
    .Y(_2673_));
 sky130_fd_sc_hd__or2_2 _5498_ (.A(_1700_),
    .B(_1703_),
    .X(_2674_));
 sky130_fd_sc_hd__nor2_4 _5499_ (.A(_2671_),
    .B(_2673_),
    .Y(_2675_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(_1469_),
    .A1(_1437_),
    .S(net194),
    .X(_2676_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_1443_),
    .B(net194),
    .Y(_2677_));
 sky130_fd_sc_hd__and3_1 _5502_ (.A(net206),
    .B(_1480_),
    .C(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__mux2_1 _5503_ (.A0(_1427_),
    .A1(_1459_),
    .S(net194),
    .X(_2679_));
 sky130_fd_sc_hd__mux2_1 _5504_ (.A0(_1488_),
    .A1(_1495_),
    .S(net194),
    .X(_2680_));
 sky130_fd_sc_hd__mux2_1 _5505_ (.A0(_2679_),
    .A1(_2680_),
    .S(net203),
    .X(_2681_));
 sky130_fd_sc_hd__a211o_1 _5506_ (.A1(net203),
    .A2(_2676_),
    .B1(_2678_),
    .C1(_1467_),
    .X(_2682_));
 sky130_fd_sc_hd__o211a_1 _5507_ (.A1(net201),
    .A2(_2681_),
    .B1(_2682_),
    .C1(net210),
    .X(_2683_));
 sky130_fd_sc_hd__mux2_1 _5508_ (.A0(_1407_),
    .A1(_1398_),
    .S(net195),
    .X(_2684_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(_1417_),
    .A1(_1381_),
    .S(net195),
    .X(_2685_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(_2684_),
    .A1(_2685_),
    .S(net203),
    .X(_2686_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(_1371_),
    .A1(_1389_),
    .S(net195),
    .X(_2687_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(_1506_),
    .A1(_1513_),
    .S(net195),
    .X(_2688_));
 sky130_fd_sc_hd__mux2_1 _5513_ (.A0(_2687_),
    .A1(_2688_),
    .S(net203),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _5514_ (.A0(_2686_),
    .A1(_2689_),
    .S(net198),
    .X(_2690_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(_1551_),
    .A1(_1559_),
    .S(net195),
    .X(_2691_));
 sky130_fd_sc_hd__mux2_1 _5516_ (.A0(_1584_),
    .A1(_1566_),
    .S(net195),
    .X(_2692_));
 sky130_fd_sc_hd__mux2_1 _5517_ (.A0(_2691_),
    .A1(_2692_),
    .S(net203),
    .X(_2693_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(_1575_),
    .A1(_1541_),
    .S(net191),
    .X(_2694_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(_1524_),
    .A1(_1533_),
    .S(net192),
    .X(_2695_));
 sky130_fd_sc_hd__mux2_1 _5520_ (.A0(_2694_),
    .A1(_2695_),
    .S(net202),
    .X(_2696_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(_2693_),
    .A1(_2696_),
    .S(net198),
    .X(_2697_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(_1648_),
    .A1(_1618_),
    .S(net191),
    .X(_2698_));
 sky130_fd_sc_hd__mux2_1 _5523_ (.A0(_1611_),
    .A1(_1627_),
    .S(net191),
    .X(_2699_));
 sky130_fd_sc_hd__mux2_1 _5524_ (.A0(_2698_),
    .A1(_2699_),
    .S(net202),
    .X(_2700_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(_1656_),
    .A1(_1603_),
    .S(net191),
    .X(_2701_));
 sky130_fd_sc_hd__mux2_1 _5526_ (.A0(_1594_),
    .A1(_1638_),
    .S(net191),
    .X(_2702_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(_2701_),
    .A1(_2702_),
    .S(net202),
    .X(_2703_));
 sky130_fd_sc_hd__mux2_2 _5528_ (.A0(_2700_),
    .A1(_2703_),
    .S(net196),
    .X(_2704_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(_2697_),
    .A1(_2704_),
    .S(net189),
    .X(_2705_));
 sky130_fd_sc_hd__a211o_1 _5530_ (.A1(net189),
    .A2(_2690_),
    .B1(_2683_),
    .C1(net214),
    .X(_2706_));
 sky130_fd_sc_hd__o21ai_1 _5531_ (.A1(net217),
    .A2(_2705_),
    .B1(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__nor3_4 _5532_ (.A(net2208),
    .B(_1700_),
    .C(_1701_),
    .Y(_2708_));
 sky130_fd_sc_hd__or3_2 _5533_ (.A(net2238),
    .B(_1700_),
    .C(_1701_),
    .X(_2709_));
 sky130_fd_sc_hd__nor2_1 _5534_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .Y(_2710_));
 sky130_fd_sc_hd__or2_4 _5535_ (.A(net2251),
    .B(net2292),
    .X(_2711_));
 sky130_fd_sc_hd__o31a_2 _5536_ (.A1(net2208),
    .A2(net2253),
    .A3(_2711_),
    .B1(net314),
    .X(_2712_));
 sky130_fd_sc_hd__nor2_8 _5537_ (.A(_1703_),
    .B(_2711_),
    .Y(_2713_));
 sky130_fd_sc_hd__or2_4 _5538_ (.A(_1703_),
    .B(_2711_),
    .X(_2714_));
 sky130_fd_sc_hd__a21o_1 _5539_ (.A1(net283),
    .A2(net312),
    .B1(_1481_),
    .X(_2715_));
 sky130_fd_sc_hd__nor2_2 _5540_ (.A(_2670_),
    .B(_2711_),
    .Y(_2716_));
 sky130_fd_sc_hd__and4bb_4 _5541_ (.A_N(net2252),
    .B_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .C(net2208),
    .D(_2710_),
    .X(_2717_));
 sky130_fd_sc_hd__nor2_8 _5542_ (.A(net310),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__or2_4 _5543_ (.A(net310),
    .B(_2717_),
    .X(_2719_));
 sky130_fd_sc_hd__nor2_8 _5544_ (.A(_1700_),
    .B(_2670_),
    .Y(_2720_));
 sky130_fd_sc_hd__or2_4 _5545_ (.A(_1700_),
    .B(_2670_),
    .X(_2721_));
 sky130_fd_sc_hd__and3_1 _5546_ (.A(_2675_),
    .B(_2718_),
    .C(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__and4_1 _5547_ (.A(_1704_),
    .B(net282),
    .C(net312),
    .D(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__nand4_4 _5548_ (.A(_1704_),
    .B(net282),
    .C(net312),
    .D(_2722_),
    .Y(_2724_));
 sky130_fd_sc_hd__a21o_1 _5549_ (.A1(net194),
    .A2(_2717_),
    .B1(net311),
    .X(_2725_));
 sky130_fd_sc_hd__a21oi_1 _5550_ (.A1(_1480_),
    .A2(_2725_),
    .B1(net221),
    .Y(_2726_));
 sky130_fd_sc_hd__nand2_4 _5551_ (.A(net217),
    .B(_2720_),
    .Y(_2727_));
 sky130_fd_sc_hd__or2_1 _5552_ (.A(net198),
    .B(_1664_),
    .X(_2728_));
 sky130_fd_sc_hd__or2_1 _5553_ (.A(net189),
    .B(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__o211a_1 _5554_ (.A1(_2727_),
    .A2(_2729_),
    .B1(_2715_),
    .C1(_2726_),
    .X(_2730_));
 sky130_fd_sc_hd__o211a_1 _5555_ (.A1(_2675_),
    .A2(_2707_),
    .B1(_2730_),
    .C1(_2669_),
    .X(_2731_));
 sky130_fd_sc_hd__a211oi_1 _5556_ (.A1(_1479_),
    .A2(net220),
    .B1(net2255),
    .C1(net460),
    .Y(_0625_));
 sky130_fd_sc_hd__mux4_1 _5557_ (.A0(_1533_),
    .A1(_1648_),
    .A2(_1541_),
    .A3(_1524_),
    .S0(net191),
    .S1(net205),
    .X(_2732_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(_1559_),
    .A1(_1584_),
    .S(net193),
    .X(_2733_));
 sky130_fd_sc_hd__mux4_1 _5559_ (.A0(_1559_),
    .A1(_1566_),
    .A2(_1584_),
    .A3(_1575_),
    .S0(net204),
    .S1(net193),
    .X(_2734_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(_2732_),
    .A1(_2734_),
    .S(net199),
    .X(_2735_));
 sky130_fd_sc_hd__nor2_1 _5561_ (.A(net186),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__mux4_1 _5562_ (.A0(_1618_),
    .A1(_1627_),
    .A2(_1611_),
    .A3(_1656_),
    .S0(net202),
    .S1(net191),
    .X(_2737_));
 sky130_fd_sc_hd__nor2_1 _5563_ (.A(net196),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__and2b_1 _5564_ (.A_N(net191),
    .B(_1603_),
    .X(_2739_));
 sky130_fd_sc_hd__a21oi_1 _5565_ (.A1(net191),
    .A2(_1594_),
    .B1(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__nand2_1 _5566_ (.A(net202),
    .B(_1638_),
    .Y(_2741_));
 sky130_fd_sc_hd__o21a_1 _5567_ (.A1(net202),
    .A2(_2740_),
    .B1(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__a21o_1 _5568_ (.A1(net196),
    .A2(_2742_),
    .B1(_2738_),
    .X(_2743_));
 sky130_fd_sc_hd__a21oi_1 _5569_ (.A1(net186),
    .A2(_2743_),
    .B1(_2736_),
    .Y(_2744_));
 sky130_fd_sc_hd__o22a_1 _5570_ (.A1(net202),
    .A2(_2740_),
    .B1(_2741_),
    .B2(net191),
    .X(_2745_));
 sky130_fd_sc_hd__a21o_1 _5571_ (.A1(net196),
    .A2(_2745_),
    .B1(_2738_),
    .X(_2746_));
 sky130_fd_sc_hd__a21oi_1 _5572_ (.A1(net187),
    .A2(_2746_),
    .B1(_2736_),
    .Y(_2747_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(net315),
    .A1(_1478_),
    .S(net194),
    .X(_2748_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(net206),
    .B(net314),
    .Y(_2749_));
 sky130_fd_sc_hd__nand2_1 _5575_ (.A(net204),
    .B(net315),
    .Y(_2750_));
 sky130_fd_sc_hd__and3_1 _5576_ (.A(_1447_),
    .B(_1448_),
    .C(net315),
    .X(_2751_));
 sky130_fd_sc_hd__a21oi_1 _5577_ (.A1(_1447_),
    .A2(_1448_),
    .B1(net315),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_1 _5578_ (.A(_2751_),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__or3_1 _5579_ (.A(_1442_),
    .B(_2751_),
    .C(_2752_),
    .X(_2754_));
 sky130_fd_sc_hd__nor2_1 _5580_ (.A(_1443_),
    .B(_2753_),
    .Y(_2755_));
 sky130_fd_sc_hd__or2_1 _5581_ (.A(_1443_),
    .B(_2753_),
    .X(_2756_));
 sky130_fd_sc_hd__nand2_1 _5582_ (.A(_2754_),
    .B(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__xor2_1 _5583_ (.A(_2748_),
    .B(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__o21a_1 _5584_ (.A1(_1443_),
    .A2(net194),
    .B1(_1479_),
    .X(_2759_));
 sky130_fd_sc_hd__inv_2 _5585_ (.A(_2759_),
    .Y(_2760_));
 sky130_fd_sc_hd__or2_1 _5586_ (.A(net203),
    .B(_2759_),
    .X(_2761_));
 sky130_fd_sc_hd__nor2_1 _5587_ (.A(net198),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__nand2_1 _5588_ (.A(net209),
    .B(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__a221oi_1 _5589_ (.A1(_1442_),
    .A2(net311),
    .B1(net281),
    .B2(net204),
    .C1(net220),
    .Y(_2764_));
 sky130_fd_sc_hd__o221a_1 _5590_ (.A1(net312),
    .A2(_2757_),
    .B1(_2763_),
    .B2(_2727_),
    .C1(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__o21ai_1 _5591_ (.A1(_2712_),
    .A2(_2758_),
    .B1(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__mux4_1 _5592_ (.A0(_1437_),
    .A1(_1442_),
    .A2(_1427_),
    .A3(_1469_),
    .S0(net206),
    .S1(net194),
    .X(_2767_));
 sky130_fd_sc_hd__mux4_2 _5593_ (.A0(_1459_),
    .A1(_1488_),
    .A2(_1495_),
    .A3(_1407_),
    .S0(_1476_),
    .S1(net204),
    .X(_2768_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(_2767_),
    .A1(_2768_),
    .S(net198),
    .X(_2769_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(_1389_),
    .A1(_1506_),
    .S(net193),
    .X(_2770_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(_1513_),
    .A1(_1551_),
    .S(net193),
    .X(_2771_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(_2770_),
    .A1(_2771_),
    .S(net204),
    .X(_2772_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(_1381_),
    .A1(_1371_),
    .S(net193),
    .X(_2773_));
 sky130_fd_sc_hd__mux4_1 _5599_ (.A0(_1381_),
    .A1(_1398_),
    .A2(_1371_),
    .A3(_1417_),
    .S0(net206),
    .S1(net193),
    .X(_2774_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(_2772_),
    .A1(_2774_),
    .S(net200),
    .X(_2775_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(_2769_),
    .A1(_2775_),
    .S(net187),
    .X(_2776_));
 sky130_fd_sc_hd__o21a_1 _5602_ (.A1(net216),
    .A2(_2747_),
    .B1(_2673_),
    .X(_2777_));
 sky130_fd_sc_hd__o21a_1 _5603_ (.A1(net216),
    .A2(_2744_),
    .B1(_2671_),
    .X(_2778_));
 sky130_fd_sc_hd__o22a_1 _5604_ (.A1(net213),
    .A2(_2776_),
    .B1(_2777_),
    .B2(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__a21o_1 _5605_ (.A1(_1442_),
    .A2(net203),
    .B1(_2724_),
    .X(_2780_));
 sky130_fd_sc_hd__o211a_1 _5606_ (.A1(_2766_),
    .A2(_2779_),
    .B1(_2780_),
    .C1(net444),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _5607_ (.A0(_2676_),
    .A1(_2679_),
    .S(net203),
    .X(_2781_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(_2680_),
    .A1(_2684_),
    .S(net203),
    .X(_2782_));
 sky130_fd_sc_hd__mux2_1 _5609_ (.A0(_2781_),
    .A1(_2782_),
    .S(net198),
    .X(_2783_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(_2685_),
    .A1(_2687_),
    .S(net203),
    .X(_2784_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(_2688_),
    .A1(_2691_),
    .S(net203),
    .X(_2785_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(_2784_),
    .A1(_2785_),
    .S(net198),
    .X(_2786_));
 sky130_fd_sc_hd__o21ba_1 _5613_ (.A1(net189),
    .A2(_2783_),
    .B1_N(_2675_),
    .X(_2787_));
 sky130_fd_sc_hd__o21ai_1 _5614_ (.A1(net210),
    .A2(_2786_),
    .B1(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__o21ai_1 _5615_ (.A1(_1469_),
    .A2(net194),
    .B1(_2677_),
    .Y(_2789_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(_1662_),
    .A1(_2789_),
    .S(net206),
    .X(_2790_));
 sky130_fd_sc_hd__or4_1 _5617_ (.A(net188),
    .B(net198),
    .C(_2721_),
    .D(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__a21oi_1 _5618_ (.A1(_2748_),
    .A2(_2754_),
    .B1(_2755_),
    .Y(_2792_));
 sky130_fd_sc_hd__a32o_1 _5619_ (.A1(_1442_),
    .A2(_2749_),
    .A3(_2750_),
    .B1(_2754_),
    .B2(_2748_),
    .X(_2793_));
 sky130_fd_sc_hd__nor2_1 _5620_ (.A(net198),
    .B(net313),
    .Y(_2794_));
 sky130_fd_sc_hd__nor2_1 _5621_ (.A(net201),
    .B(net315),
    .Y(_2795_));
 sky130_fd_sc_hd__or3_1 _5622_ (.A(_1469_),
    .B(_2794_),
    .C(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__o21ai_1 _5623_ (.A1(_2794_),
    .A2(_2795_),
    .B1(_1469_),
    .Y(_2797_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(_2796_),
    .B(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__a21oi_1 _5625_ (.A1(_2792_),
    .A2(_2798_),
    .B1(net283),
    .Y(_2799_));
 sky130_fd_sc_hd__o21a_1 _5626_ (.A1(_2792_),
    .A2(_2798_),
    .B1(_2799_),
    .X(_2800_));
 sky130_fd_sc_hd__a221o_1 _5627_ (.A1(_1469_),
    .A2(_2716_),
    .B1(net281),
    .B2(net198),
    .C1(net221),
    .X(_2801_));
 sky130_fd_sc_hd__nor2_1 _5628_ (.A(_1470_),
    .B(net312),
    .Y(_2802_));
 sky130_fd_sc_hd__mux2_1 _5629_ (.A0(_2692_),
    .A1(_2694_),
    .S(net203),
    .X(_2803_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(_2695_),
    .A1(_2698_),
    .S(net202),
    .X(_2804_));
 sky130_fd_sc_hd__mux2_1 _5631_ (.A0(_2803_),
    .A1(_2804_),
    .S(net197),
    .X(_2805_));
 sky130_fd_sc_hd__nor2_1 _5632_ (.A(net188),
    .B(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(_2699_),
    .A1(_2701_),
    .S(net202),
    .X(_2807_));
 sky130_fd_sc_hd__nor2_1 _5634_ (.A(net196),
    .B(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(net205),
    .B(_2702_),
    .Y(_2809_));
 sky130_fd_sc_hd__and2_1 _5636_ (.A(_2741_),
    .B(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__a21oi_1 _5637_ (.A1(net196),
    .A2(_2810_),
    .B1(_2808_),
    .Y(_2811_));
 sky130_fd_sc_hd__nor2_1 _5638_ (.A(net207),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__a21oi_1 _5639_ (.A1(net196),
    .A2(_2809_),
    .B1(_2808_),
    .Y(_2813_));
 sky130_fd_sc_hd__inv_2 _5640_ (.A(_2813_),
    .Y(_2814_));
 sky130_fd_sc_hd__a211o_1 _5641_ (.A1(net186),
    .A2(_2814_),
    .B1(_2806_),
    .C1(_2674_),
    .X(_2815_));
 sky130_fd_sc_hd__o311a_1 _5642_ (.A1(_2672_),
    .A2(_2806_),
    .A3(_2812_),
    .B1(_2815_),
    .C1(net212),
    .X(_2816_));
 sky130_fd_sc_hd__a31o_1 _5643_ (.A1(net217),
    .A2(_2788_),
    .A3(_2791_),
    .B1(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__or4b_1 _5644_ (.A(_2800_),
    .B(_2801_),
    .C(_2802_),
    .D_N(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__a21o_1 _5645_ (.A1(net198),
    .A2(_1469_),
    .B1(net219),
    .X(_2819_));
 sky130_fd_sc_hd__and3_1 _5646_ (.A(net444),
    .B(_2818_),
    .C(net2338),
    .X(_0627_));
 sky130_fd_sc_hd__mux4_1 _5647_ (.A0(_1541_),
    .A1(_1566_),
    .A2(_1524_),
    .A3(_1575_),
    .S0(net205),
    .S1(net192),
    .X(_2820_));
 sky130_fd_sc_hd__mux4_1 _5648_ (.A0(_1533_),
    .A1(_1618_),
    .A2(_1648_),
    .A3(_1611_),
    .S0(net202),
    .S1(net192),
    .X(_2821_));
 sky130_fd_sc_hd__mux2_1 _5649_ (.A0(_2820_),
    .A1(_2821_),
    .S(net197),
    .X(_2822_));
 sky130_fd_sc_hd__nor2_1 _5650_ (.A(net186),
    .B(_2822_),
    .Y(_2823_));
 sky130_fd_sc_hd__mux4_1 _5651_ (.A0(_1603_),
    .A1(_1627_),
    .A2(_1594_),
    .A3(_1656_),
    .S0(net205),
    .S1(net191),
    .X(_2824_));
 sky130_fd_sc_hd__and2_1 _5652_ (.A(net199),
    .B(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__nor2_1 _5653_ (.A(net199),
    .B(net190),
    .Y(_2826_));
 sky130_fd_sc_hd__nand2_1 _5654_ (.A(net196),
    .B(_1638_),
    .Y(_2827_));
 sky130_fd_sc_hd__nor2_1 _5655_ (.A(_2825_),
    .B(_2826_),
    .Y(_2828_));
 sky130_fd_sc_hd__a21oi_1 _5656_ (.A1(net186),
    .A2(_2828_),
    .B1(_2823_),
    .Y(_2829_));
 sky130_fd_sc_hd__nor3_1 _5657_ (.A(net202),
    .B(net192),
    .C(net190),
    .Y(_2830_));
 sky130_fd_sc_hd__a21oi_1 _5658_ (.A1(net197),
    .A2(_2830_),
    .B1(_2825_),
    .Y(_2831_));
 sky130_fd_sc_hd__a21oi_1 _5659_ (.A1(net186),
    .A2(_2831_),
    .B1(_2823_),
    .Y(_2832_));
 sky130_fd_sc_hd__a21bo_1 _5660_ (.A1(_2793_),
    .A2(_2796_),
    .B1_N(_2797_),
    .X(_2833_));
 sky130_fd_sc_hd__xnor2_1 _5661_ (.A(net210),
    .B(net315),
    .Y(_2834_));
 sky130_fd_sc_hd__or2_1 _5662_ (.A(_1437_),
    .B(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__nand2_1 _5663_ (.A(_1437_),
    .B(_2834_),
    .Y(_2836_));
 sky130_fd_sc_hd__nand2_1 _5664_ (.A(_2835_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__xor2_1 _5665_ (.A(_2833_),
    .B(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__a21oi_1 _5666_ (.A1(_1437_),
    .A2(net311),
    .B1(net189),
    .Y(_2839_));
 sky130_fd_sc_hd__o221a_1 _5667_ (.A1(_2714_),
    .A2(_2837_),
    .B1(_2839_),
    .B2(_2718_),
    .C1(net219),
    .X(_2840_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(_1437_),
    .A1(_1469_),
    .S(net194),
    .X(_2841_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(_2760_),
    .A1(_2841_),
    .S(_1449_),
    .X(_2842_));
 sky130_fd_sc_hd__nand2_1 _5670_ (.A(net201),
    .B(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__o31a_1 _5671_ (.A1(net189),
    .A2(_2727_),
    .A3(_2843_),
    .B1(_2840_),
    .X(_2844_));
 sky130_fd_sc_hd__mux4_1 _5672_ (.A0(_1437_),
    .A1(_1459_),
    .A2(_1427_),
    .A3(_1488_),
    .S0(net203),
    .S1(net194),
    .X(_2845_));
 sky130_fd_sc_hd__mux4_1 _5673_ (.A0(_1398_),
    .A1(_1417_),
    .A2(_1495_),
    .A3(_1407_),
    .S0(net195),
    .S1(net206),
    .X(_2846_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(_2845_),
    .A1(_2846_),
    .S(net198),
    .X(_2847_));
 sky130_fd_sc_hd__mux2_1 _5675_ (.A0(_2770_),
    .A1(_2773_),
    .S(net206),
    .X(_2848_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(_2733_),
    .A1(_2771_),
    .S(net205),
    .X(_2849_));
 sky130_fd_sc_hd__mux2_1 _5677_ (.A0(_2848_),
    .A1(_2849_),
    .S(net197),
    .X(_2850_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(_2847_),
    .A1(_2850_),
    .S(net186),
    .X(_2851_));
 sky130_fd_sc_hd__o21a_1 _5679_ (.A1(net215),
    .A2(_2832_),
    .B1(_2673_),
    .X(_2852_));
 sky130_fd_sc_hd__o21a_1 _5680_ (.A1(net215),
    .A2(_2829_),
    .B1(_2671_),
    .X(_2853_));
 sky130_fd_sc_hd__o22a_2 _5681_ (.A1(net212),
    .A2(_2851_),
    .B1(_2852_),
    .B2(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__o21ai_1 _5682_ (.A1(net283),
    .A2(_2838_),
    .B1(_2844_),
    .Y(_2855_));
 sky130_fd_sc_hd__a21o_1 _5683_ (.A1(net189),
    .A2(_1437_),
    .B1(net219),
    .X(_2856_));
 sky130_fd_sc_hd__o211a_1 _5684_ (.A1(_2854_),
    .A2(_2855_),
    .B1(_2856_),
    .C1(net444),
    .X(_0628_));
 sky130_fd_sc_hd__a21bo_1 _5685_ (.A1(_2833_),
    .A2(_2835_),
    .B1_N(_2836_),
    .X(_2857_));
 sky130_fd_sc_hd__xnor2_1 _5686_ (.A(net217),
    .B(net315),
    .Y(_2858_));
 sky130_fd_sc_hd__nor2_1 _5687_ (.A(_1427_),
    .B(_2858_),
    .Y(_2859_));
 sky130_fd_sc_hd__or2_1 _5688_ (.A(_1427_),
    .B(_2858_),
    .X(_2860_));
 sky130_fd_sc_hd__and2_1 _5689_ (.A(_1427_),
    .B(_2858_),
    .X(_2861_));
 sky130_fd_sc_hd__nor2_1 _5690_ (.A(_2859_),
    .B(_2861_),
    .Y(_2862_));
 sky130_fd_sc_hd__a21oi_1 _5691_ (.A1(_2857_),
    .A2(_2862_),
    .B1(net283),
    .Y(_2863_));
 sky130_fd_sc_hd__o21ai_1 _5692_ (.A1(_2857_),
    .A2(_2862_),
    .B1(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(_2696_),
    .A1(_2700_),
    .S(net196),
    .X(_2865_));
 sky130_fd_sc_hd__nand2_1 _5694_ (.A(net208),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__and2_1 _5695_ (.A(net199),
    .B(_2703_),
    .X(_2867_));
 sky130_fd_sc_hd__nor2_1 _5696_ (.A(_2826_),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__o21ai_1 _5697_ (.A1(net208),
    .A2(_2868_),
    .B1(_2866_),
    .Y(_2869_));
 sky130_fd_sc_hd__o311a_1 _5698_ (.A1(net208),
    .A2(_2671_),
    .A3(_2867_),
    .B1(_2869_),
    .C1(net212),
    .X(_2870_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(_2689_),
    .A1(_2693_),
    .S(net198),
    .X(_2871_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(_2681_),
    .A1(_2686_),
    .S(net198),
    .X(_2872_));
 sky130_fd_sc_hd__or2_1 _5701_ (.A(net189),
    .B(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__o211a_1 _5702_ (.A1(net210),
    .A2(_2871_),
    .B1(_2873_),
    .C1(net217),
    .X(_2874_));
 sky130_fd_sc_hd__nor2_1 _5703_ (.A(_2870_),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__a221o_1 _5704_ (.A1(_1428_),
    .A2(_2713_),
    .B1(_2717_),
    .B2(net214),
    .C1(net311),
    .X(_2876_));
 sky130_fd_sc_hd__a21oi_1 _5705_ (.A1(_1429_),
    .A2(_2876_),
    .B1(net221),
    .Y(_2877_));
 sky130_fd_sc_hd__mux4_1 _5706_ (.A0(_1427_),
    .A1(_1437_),
    .A2(_1469_),
    .A3(_1442_),
    .S0(net194),
    .S1(net204),
    .X(_2878_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(_1665_),
    .A1(_2878_),
    .S(net201),
    .X(_2879_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(net210),
    .B(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__o221a_1 _5709_ (.A1(_2675_),
    .A2(_2875_),
    .B1(_2880_),
    .B2(_2727_),
    .C1(_2877_),
    .X(_2881_));
 sky130_fd_sc_hd__a221oi_1 _5710_ (.A1(_1428_),
    .A2(net221),
    .B1(_2864_),
    .B2(_2881_),
    .C1(net460),
    .Y(_0629_));
 sky130_fd_sc_hd__xnor2_1 _5711_ (.A(_1457_),
    .B(net314),
    .Y(_2882_));
 sky130_fd_sc_hd__nor2_1 _5712_ (.A(_1459_),
    .B(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__nand2_1 _5713_ (.A(_1459_),
    .B(_2882_),
    .Y(_2884_));
 sky130_fd_sc_hd__nand2b_1 _5714_ (.A_N(_2883_),
    .B(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__a21oi_2 _5715_ (.A1(_2857_),
    .A2(_2860_),
    .B1(_2861_),
    .Y(_2886_));
 sky130_fd_sc_hd__xnor2_1 _5716_ (.A(_2885_),
    .B(_2886_),
    .Y(_2887_));
 sky130_fd_sc_hd__nor2_1 _5717_ (.A(net283),
    .B(_2887_),
    .Y(_2888_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(_2732_),
    .A1(_2737_),
    .S(net196),
    .X(_2889_));
 sky130_fd_sc_hd__nor2_1 _5719_ (.A(net187),
    .B(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__nor2_1 _5720_ (.A(net196),
    .B(_2745_),
    .Y(_2891_));
 sky130_fd_sc_hd__inv_2 _5721_ (.A(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__a211o_1 _5722_ (.A1(net187),
    .A2(_2892_),
    .B1(_2890_),
    .C1(_2674_),
    .X(_2893_));
 sky130_fd_sc_hd__o21a_1 _5723_ (.A1(net196),
    .A2(_2742_),
    .B1(_2827_),
    .X(_2894_));
 sky130_fd_sc_hd__a21oi_1 _5724_ (.A1(net187),
    .A2(_2894_),
    .B1(_2890_),
    .Y(_2895_));
 sky130_fd_sc_hd__a21bo_2 _5725_ (.A1(_2671_),
    .A2(_2895_),
    .B1_N(_2893_),
    .X(_2896_));
 sky130_fd_sc_hd__a221o_1 _5726_ (.A1(_1459_),
    .A2(net311),
    .B1(net281),
    .B2(_1457_),
    .C1(net221),
    .X(_2897_));
 sky130_fd_sc_hd__nor2_1 _5727_ (.A(net312),
    .B(_2885_),
    .Y(_2898_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(_1459_),
    .A1(_1427_),
    .S(net194),
    .X(_2899_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(_2841_),
    .A1(_2899_),
    .S(_1449_),
    .X(_2900_));
 sky130_fd_sc_hd__inv_2 _5730_ (.A(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__mux2_1 _5731_ (.A0(_2761_),
    .A1(_2901_),
    .S(net200),
    .X(_2902_));
 sky130_fd_sc_hd__or3_2 _5732_ (.A(net188),
    .B(_2721_),
    .C(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_1 _5733_ (.A0(_2768_),
    .A1(_2774_),
    .S(net197),
    .X(_2904_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(_2734_),
    .A1(_2772_),
    .S(net200),
    .X(_2905_));
 sky130_fd_sc_hd__o21ba_1 _5735_ (.A1(net209),
    .A2(_2905_),
    .B1_N(_2675_),
    .X(_2906_));
 sky130_fd_sc_hd__o21ai_2 _5736_ (.A1(net186),
    .A2(_2904_),
    .B1(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__a21oi_4 _5737_ (.A1(_2903_),
    .A2(_2907_),
    .B1(net213),
    .Y(_2908_));
 sky130_fd_sc_hd__a211o_1 _5738_ (.A1(net214),
    .A2(_2896_),
    .B1(_2897_),
    .C1(_2898_),
    .X(_2909_));
 sky130_fd_sc_hd__a21o_1 _5739_ (.A1(_1457_),
    .A2(_1459_),
    .B1(net219),
    .X(_2910_));
 sky130_fd_sc_hd__o311a_2 _5740_ (.A1(_2888_),
    .A2(_2908_),
    .A3(_2909_),
    .B1(net2312),
    .C1(net444),
    .X(_0630_));
 sky130_fd_sc_hd__o21ai_2 _5741_ (.A1(_2883_),
    .A2(_2886_),
    .B1(_2884_),
    .Y(_2911_));
 sky130_fd_sc_hd__xnor2_1 _5742_ (.A(_1486_),
    .B(net313),
    .Y(_2912_));
 sky130_fd_sc_hd__nor2_1 _5743_ (.A(_1488_),
    .B(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__or2_1 _5744_ (.A(_1488_),
    .B(_2912_),
    .X(_2914_));
 sky130_fd_sc_hd__and2_1 _5745_ (.A(_1488_),
    .B(_2912_),
    .X(_2915_));
 sky130_fd_sc_hd__nor2_1 _5746_ (.A(_2913_),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__a21oi_1 _5747_ (.A1(_2911_),
    .A2(_2916_),
    .B1(net283),
    .Y(_2917_));
 sky130_fd_sc_hd__o21a_1 _5748_ (.A1(_2911_),
    .A2(_2916_),
    .B1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(_2804_),
    .A1(_2807_),
    .S(net196),
    .X(_2919_));
 sky130_fd_sc_hd__or2_1 _5750_ (.A(net187),
    .B(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__nor2_1 _5751_ (.A(net187),
    .B(_2674_),
    .Y(_2921_));
 sky130_fd_sc_hd__nand2_2 _5752_ (.A(net207),
    .B(_2673_),
    .Y(_2922_));
 sky130_fd_sc_hd__or2_1 _5753_ (.A(net196),
    .B(_2809_),
    .X(_2923_));
 sky130_fd_sc_hd__nor2_1 _5754_ (.A(_2674_),
    .B(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__o21a_1 _5755_ (.A1(_2921_),
    .A2(_2924_),
    .B1(_2920_),
    .X(_2925_));
 sky130_fd_sc_hd__o21ai_2 _5756_ (.A1(net196),
    .A2(_2810_),
    .B1(_2827_),
    .Y(_2926_));
 sky130_fd_sc_hd__o211a_1 _5757_ (.A1(net207),
    .A2(_2926_),
    .B1(_2920_),
    .C1(_2671_),
    .X(_2927_));
 sky130_fd_sc_hd__o21ai_1 _5758_ (.A1(_2925_),
    .A2(_2927_),
    .B1(net211),
    .Y(_2928_));
 sky130_fd_sc_hd__a21o_1 _5759_ (.A1(_1488_),
    .A2(net311),
    .B1(_1486_),
    .X(_2929_));
 sky130_fd_sc_hd__a221o_1 _5760_ (.A1(_1489_),
    .A2(_2713_),
    .B1(net281),
    .B2(_2929_),
    .C1(net220),
    .X(_2930_));
 sky130_fd_sc_hd__mux4_2 _5761_ (.A0(_1427_),
    .A1(_1437_),
    .A2(_1488_),
    .A3(_1459_),
    .S0(_1476_),
    .S1(net206),
    .X(_2931_));
 sky130_fd_sc_hd__inv_2 _5762_ (.A(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(_2790_),
    .A1(_2932_),
    .S(net200),
    .X(_2933_));
 sky130_fd_sc_hd__or3_2 _5764_ (.A(net188),
    .B(_2721_),
    .C(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(_2782_),
    .A1(_2784_),
    .S(net198),
    .X(_2935_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(_2785_),
    .A1(_2803_),
    .S(net198),
    .X(_2936_));
 sky130_fd_sc_hd__nor2_1 _5767_ (.A(net189),
    .B(_2935_),
    .Y(_2937_));
 sky130_fd_sc_hd__nor2_1 _5768_ (.A(net210),
    .B(_2936_),
    .Y(_2938_));
 sky130_fd_sc_hd__o31a_1 _5769_ (.A1(_2675_),
    .A2(_2937_),
    .A3(_2938_),
    .B1(_2934_),
    .X(_2939_));
 sky130_fd_sc_hd__o21ai_1 _5770_ (.A1(net214),
    .A2(_2939_),
    .B1(_2928_),
    .Y(_2940_));
 sky130_fd_sc_hd__a21o_1 _5771_ (.A1(_1486_),
    .A2(net2266),
    .B1(net219),
    .X(_2941_));
 sky130_fd_sc_hd__o311a_1 _5772_ (.A1(_2918_),
    .A2(_2930_),
    .A3(_2940_),
    .B1(_2941_),
    .C1(net444),
    .X(_0631_));
 sky130_fd_sc_hd__xnor2_1 _5773_ (.A(_1493_),
    .B(net313),
    .Y(_2942_));
 sky130_fd_sc_hd__or2_1 _5774_ (.A(_1495_),
    .B(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__nand2_1 _5775_ (.A(_1495_),
    .B(_2942_),
    .Y(_2944_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_2943_),
    .B(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__a21o_1 _5777_ (.A1(_2911_),
    .A2(_2914_),
    .B1(_2915_),
    .X(_2946_));
 sky130_fd_sc_hd__nand2_1 _5778_ (.A(_2945_),
    .B(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__or2_1 _5779_ (.A(_2945_),
    .B(_2946_),
    .X(_2948_));
 sky130_fd_sc_hd__a21oi_1 _5780_ (.A1(_2947_),
    .A2(_2948_),
    .B1(net283),
    .Y(_2949_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(_1495_),
    .A1(_1488_),
    .S(net195),
    .X(_2950_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(_2899_),
    .A1(_2950_),
    .S(net206),
    .X(_2951_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(_2842_),
    .A1(_2951_),
    .S(net200),
    .X(_2952_));
 sky130_fd_sc_hd__or3b_2 _5784_ (.A(net188),
    .B(_2721_),
    .C_N(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(_2846_),
    .A1(_2848_),
    .S(net197),
    .X(_2954_));
 sky130_fd_sc_hd__mux2_1 _5786_ (.A0(_2820_),
    .A1(_2849_),
    .S(net200),
    .X(_2955_));
 sky130_fd_sc_hd__nor2_1 _5787_ (.A(net188),
    .B(_2954_),
    .Y(_2956_));
 sky130_fd_sc_hd__nor2_1 _5788_ (.A(net210),
    .B(_2955_),
    .Y(_2957_));
 sky130_fd_sc_hd__o31a_2 _5789_ (.A1(_2675_),
    .A2(_2956_),
    .A3(_2957_),
    .B1(_2953_),
    .X(_2958_));
 sky130_fd_sc_hd__a221o_1 _5790_ (.A1(_1495_),
    .A2(net311),
    .B1(_2719_),
    .B2(_1493_),
    .C1(net221),
    .X(_2959_));
 sky130_fd_sc_hd__o22ai_1 _5791_ (.A1(_2714_),
    .A2(_2945_),
    .B1(_2958_),
    .B2(_1425_),
    .Y(_2960_));
 sky130_fd_sc_hd__mux2_1 _5792_ (.A0(_2821_),
    .A1(_2824_),
    .S(net197),
    .X(_2961_));
 sky130_fd_sc_hd__or2_1 _5793_ (.A(net187),
    .B(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__a21o_1 _5794_ (.A1(net199),
    .A2(_2830_),
    .B1(net208),
    .X(_2963_));
 sky130_fd_sc_hd__and3_1 _5795_ (.A(_2673_),
    .B(_2962_),
    .C(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__o21a_1 _5796_ (.A1(net207),
    .A2(_1638_),
    .B1(_2962_),
    .X(_2965_));
 sky130_fd_sc_hd__a21o_2 _5797_ (.A1(_2671_),
    .A2(_2965_),
    .B1(_2964_),
    .X(_2966_));
 sky130_fd_sc_hd__a211o_1 _5798_ (.A1(_1425_),
    .A2(_2966_),
    .B1(_2960_),
    .C1(_2959_),
    .X(_2967_));
 sky130_fd_sc_hd__a21o_1 _5799_ (.A1(_1493_),
    .A2(_1495_),
    .B1(_2724_),
    .X(_2968_));
 sky130_fd_sc_hd__o211a_1 _5800_ (.A1(_2949_),
    .A2(_2967_),
    .B1(_2968_),
    .C1(net444),
    .X(_0632_));
 sky130_fd_sc_hd__a21bo_1 _5801_ (.A1(_2943_),
    .A2(_2946_),
    .B1_N(_2944_),
    .X(_2969_));
 sky130_fd_sc_hd__xnor2_1 _5802_ (.A(_1405_),
    .B(net314),
    .Y(_2970_));
 sky130_fd_sc_hd__nor2_1 _5803_ (.A(_1407_),
    .B(_2970_),
    .Y(_2971_));
 sky130_fd_sc_hd__or2_1 _5804_ (.A(_1407_),
    .B(_2970_),
    .X(_2972_));
 sky130_fd_sc_hd__and2_1 _5805_ (.A(_1407_),
    .B(_2970_),
    .X(_2973_));
 sky130_fd_sc_hd__nor2_1 _5806_ (.A(_2971_),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__xnor2_1 _5807_ (.A(_2969_),
    .B(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__a21o_1 _5808_ (.A1(_1407_),
    .A2(net311),
    .B1(_1405_),
    .X(_2976_));
 sky130_fd_sc_hd__a221o_1 _5809_ (.A1(_1410_),
    .A2(_2713_),
    .B1(_2719_),
    .B2(_2976_),
    .C1(net221),
    .X(_2977_));
 sky130_fd_sc_hd__mux4_1 _5810_ (.A0(_1407_),
    .A1(_1488_),
    .A2(_1495_),
    .A3(_1459_),
    .S0(net203),
    .S1(net194),
    .X(_2978_));
 sky130_fd_sc_hd__mux2_1 _5811_ (.A0(_2878_),
    .A1(_2978_),
    .S(net201),
    .X(_2979_));
 sky130_fd_sc_hd__inv_2 _5812_ (.A(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__mux2_1 _5813_ (.A0(_2728_),
    .A1(_2980_),
    .S(net210),
    .X(_2981_));
 sky130_fd_sc_hd__mux2_1 _5814_ (.A0(_2690_),
    .A1(_2697_),
    .S(net189),
    .X(_2982_));
 sky130_fd_sc_hd__nor2_1 _5815_ (.A(net214),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__o22a_1 _5816_ (.A1(_2721_),
    .A2(_2981_),
    .B1(_2983_),
    .B2(_2675_),
    .X(_2984_));
 sky130_fd_sc_hd__nand2_1 _5817_ (.A(net207),
    .B(_2704_),
    .Y(_2985_));
 sky130_fd_sc_hd__or2_2 _5818_ (.A(net207),
    .B(net190),
    .X(_2986_));
 sky130_fd_sc_hd__o221a_1 _5819_ (.A1(_2675_),
    .A2(_2985_),
    .B1(_2986_),
    .B2(_2672_),
    .C1(net212),
    .X(_2987_));
 sky130_fd_sc_hd__o22ai_1 _5820_ (.A1(net283),
    .A2(_2975_),
    .B1(_2984_),
    .B2(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__a21o_1 _5821_ (.A1(_1405_),
    .A2(_1407_),
    .B1(net219),
    .X(_2989_));
 sky130_fd_sc_hd__o211a_1 _5822_ (.A1(_2977_),
    .A2(_2988_),
    .B1(_2989_),
    .C1(net444),
    .X(_0633_));
 sky130_fd_sc_hd__xnor2_1 _5823_ (.A(_1396_),
    .B(net313),
    .Y(_2990_));
 sky130_fd_sc_hd__or2_1 _5824_ (.A(_1398_),
    .B(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__and2_1 _5825_ (.A(_1398_),
    .B(_2990_),
    .X(_2992_));
 sky130_fd_sc_hd__inv_2 _5826_ (.A(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_2991_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__a21o_1 _5828_ (.A1(_2969_),
    .A2(_2972_),
    .B1(_2973_),
    .X(_2995_));
 sky130_fd_sc_hd__xor2_1 _5829_ (.A(_2994_),
    .B(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(_1398_),
    .A1(_1407_),
    .S(net195),
    .X(_2997_));
 sky130_fd_sc_hd__mux2_1 _5831_ (.A0(_2950_),
    .A1(_2997_),
    .S(net206),
    .X(_2998_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(_2900_),
    .A1(_2998_),
    .S(net200),
    .X(_2999_));
 sky130_fd_sc_hd__mux2_1 _5833_ (.A0(_2762_),
    .A1(_2999_),
    .S(net209),
    .X(_3000_));
 sky130_fd_sc_hd__mux2_1 _5834_ (.A0(_2735_),
    .A1(_2775_),
    .S(net209),
    .X(_3001_));
 sky130_fd_sc_hd__inv_2 _5835_ (.A(_3001_),
    .Y(_3002_));
 sky130_fd_sc_hd__o2bb2a_1 _5836_ (.A1_N(_2720_),
    .A2_N(_3000_),
    .B1(_3002_),
    .B2(_2675_),
    .X(_3003_));
 sky130_fd_sc_hd__a21oi_1 _5837_ (.A1(_1398_),
    .A2(net311),
    .B1(_1396_),
    .Y(_3004_));
 sky130_fd_sc_hd__o221a_1 _5838_ (.A1(net312),
    .A2(_2994_),
    .B1(_3004_),
    .B2(_2718_),
    .C1(net218),
    .X(_3005_));
 sky130_fd_sc_hd__mux2_1 _5839_ (.A0(_1637_),
    .A1(_2743_),
    .S(net207),
    .X(_3006_));
 sky130_fd_sc_hd__o22a_1 _5840_ (.A1(_2746_),
    .A2(_2922_),
    .B1(_3006_),
    .B2(_2672_),
    .X(_3007_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(_3003_),
    .A1(_3007_),
    .S(net213),
    .X(_3008_));
 sky130_fd_sc_hd__o211a_1 _5842_ (.A1(net283),
    .A2(_2996_),
    .B1(_3005_),
    .C1(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__a21oi_1 _5843_ (.A1(net2303),
    .A2(_1398_),
    .B1(net218),
    .Y(_3010_));
 sky130_fd_sc_hd__nor3_1 _5844_ (.A(net63),
    .B(_3009_),
    .C(net2304),
    .Y(_0634_));
 sky130_fd_sc_hd__a21oi_2 _5845_ (.A1(_2991_),
    .A2(_2995_),
    .B1(_2992_),
    .Y(_3011_));
 sky130_fd_sc_hd__xnor2_1 _5846_ (.A(_1415_),
    .B(net313),
    .Y(_3012_));
 sky130_fd_sc_hd__nor2_1 _5847_ (.A(_1417_),
    .B(_3012_),
    .Y(_3013_));
 sky130_fd_sc_hd__nand2_1 _5848_ (.A(_1417_),
    .B(_3012_),
    .Y(_3014_));
 sky130_fd_sc_hd__nand2b_1 _5849_ (.A_N(_3013_),
    .B(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__xnor2_1 _5850_ (.A(_3011_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__nor2_1 _5851_ (.A(net283),
    .B(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_2813_),
    .B(_2921_),
    .Y(_3018_));
 sky130_fd_sc_hd__a21boi_1 _5853_ (.A1(net207),
    .A2(_2811_),
    .B1_N(_2986_),
    .Y(_3019_));
 sky130_fd_sc_hd__o21ai_1 _5854_ (.A1(_2672_),
    .A2(_3019_),
    .B1(_3018_),
    .Y(_3020_));
 sky130_fd_sc_hd__a221o_1 _5855_ (.A1(_1417_),
    .A2(net310),
    .B1(net281),
    .B2(_1415_),
    .C1(net220),
    .X(_3021_));
 sky130_fd_sc_hd__nor2_1 _5856_ (.A(_1418_),
    .B(_2714_),
    .Y(_3022_));
 sky130_fd_sc_hd__a211o_1 _5857_ (.A1(net212),
    .A2(_3020_),
    .B1(_3021_),
    .C1(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__mux4_1 _5858_ (.A0(_1407_),
    .A1(_1495_),
    .A2(_1417_),
    .A3(_1398_),
    .S0(net195),
    .S1(net206),
    .X(_3024_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(_2931_),
    .A1(_3024_),
    .S(net200),
    .X(_3025_));
 sky130_fd_sc_hd__o21ai_1 _5860_ (.A1(net197),
    .A2(_2790_),
    .B1(net188),
    .Y(_3026_));
 sky130_fd_sc_hd__o211ai_2 _5861_ (.A1(net188),
    .A2(_3025_),
    .B1(_3026_),
    .C1(_2720_),
    .Y(_3027_));
 sky130_fd_sc_hd__o21ba_1 _5862_ (.A1(net188),
    .A2(_2786_),
    .B1_N(_2675_),
    .X(_3028_));
 sky130_fd_sc_hd__o21ai_1 _5863_ (.A1(net209),
    .A2(_2805_),
    .B1(_3028_),
    .Y(_3029_));
 sky130_fd_sc_hd__a21oi_1 _5864_ (.A1(_3027_),
    .A2(_3029_),
    .B1(net213),
    .Y(_3030_));
 sky130_fd_sc_hd__a21o_1 _5865_ (.A1(_1415_),
    .A2(_1417_),
    .B1(net219),
    .X(_3031_));
 sky130_fd_sc_hd__o311a_1 _5866_ (.A1(_3017_),
    .A2(_3023_),
    .A3(_3030_),
    .B1(_3031_),
    .C1(net440),
    .X(_0635_));
 sky130_fd_sc_hd__xnor2_1 _5867_ (.A(_1378_),
    .B(net316),
    .Y(_3032_));
 sky130_fd_sc_hd__or2_1 _5868_ (.A(_1381_),
    .B(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__and2_1 _5869_ (.A(_1381_),
    .B(_3032_),
    .X(_3034_));
 sky130_fd_sc_hd__inv_2 _5870_ (.A(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_3033_),
    .B(_3035_),
    .Y(_3036_));
 sky130_fd_sc_hd__o21ai_2 _5872_ (.A1(_3011_),
    .A2(_3013_),
    .B1(_3014_),
    .Y(_3037_));
 sky130_fd_sc_hd__xor2_1 _5873_ (.A(_3036_),
    .B(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__a21oi_1 _5874_ (.A1(_1381_),
    .A2(net310),
    .B1(_1379_),
    .Y(_3039_));
 sky130_fd_sc_hd__o221a_1 _5875_ (.A1(net312),
    .A2(_3036_),
    .B1(_3039_),
    .B2(_2718_),
    .C1(net218),
    .X(_3040_));
 sky130_fd_sc_hd__o21a_1 _5876_ (.A1(net187),
    .A2(_2828_),
    .B1(_2986_),
    .X(_3041_));
 sky130_fd_sc_hd__o221a_1 _5877_ (.A1(_2831_),
    .A2(_2922_),
    .B1(_3041_),
    .B2(_2672_),
    .C1(net211),
    .X(_3042_));
 sky130_fd_sc_hd__o21ba_1 _5878_ (.A1(net186),
    .A2(_2850_),
    .B1_N(_2675_),
    .X(_3043_));
 sky130_fd_sc_hd__o21ai_1 _5879_ (.A1(net208),
    .A2(_2822_),
    .B1(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(_1381_),
    .A1(_1417_),
    .S(net195),
    .X(_3045_));
 sky130_fd_sc_hd__mux2_1 _5881_ (.A0(_2997_),
    .A1(_3045_),
    .S(_1449_),
    .X(_3046_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(_2951_),
    .A1(_3046_),
    .S(net200),
    .X(_3047_));
 sky130_fd_sc_hd__nor2_1 _5883_ (.A(net188),
    .B(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__a211o_1 _5884_ (.A1(net188),
    .A2(_2843_),
    .B1(_3048_),
    .C1(_2721_),
    .X(_3049_));
 sky130_fd_sc_hd__a31o_1 _5885_ (.A1(net215),
    .A2(_3044_),
    .A3(_3049_),
    .B1(_3042_),
    .X(_3050_));
 sky130_fd_sc_hd__o211ai_1 _5886_ (.A1(net282),
    .A2(_3038_),
    .B1(_3040_),
    .C1(_3050_),
    .Y(_3051_));
 sky130_fd_sc_hd__a21o_1 _5887_ (.A1(_1379_),
    .A2(_1381_),
    .B1(net218),
    .X(_3052_));
 sky130_fd_sc_hd__and3_1 _5888_ (.A(net435),
    .B(_3051_),
    .C(_3052_),
    .X(_0636_));
 sky130_fd_sc_hd__a21oi_2 _5889_ (.A1(_3033_),
    .A2(_3037_),
    .B1(_3034_),
    .Y(_3053_));
 sky130_fd_sc_hd__xnor2_1 _5890_ (.A(_1354_),
    .B(net313),
    .Y(_3054_));
 sky130_fd_sc_hd__nor2_1 _5891_ (.A(_1371_),
    .B(_3054_),
    .Y(_3055_));
 sky130_fd_sc_hd__nand2_1 _5892_ (.A(_1371_),
    .B(_3054_),
    .Y(_3056_));
 sky130_fd_sc_hd__nand2b_1 _5893_ (.A_N(_3055_),
    .B(_3056_),
    .Y(_3057_));
 sky130_fd_sc_hd__xnor2_1 _5894_ (.A(_3053_),
    .B(_3057_),
    .Y(_3058_));
 sky130_fd_sc_hd__o21a_1 _5895_ (.A1(net187),
    .A2(_2868_),
    .B1(_2986_),
    .X(_3059_));
 sky130_fd_sc_hd__a2bb2o_1 _5896_ (.A1_N(_2672_),
    .A2_N(_3059_),
    .B1(_2921_),
    .B2(_2867_),
    .X(_3060_));
 sky130_fd_sc_hd__a221o_1 _5897_ (.A1(_1371_),
    .A2(net311),
    .B1(net281),
    .B2(_1354_),
    .C1(net220),
    .X(_3061_));
 sky130_fd_sc_hd__a22o_1 _5898_ (.A1(_1373_),
    .A2(_2713_),
    .B1(_3060_),
    .B2(net211),
    .X(_3062_));
 sky130_fd_sc_hd__mux4_1 _5899_ (.A0(_1371_),
    .A1(_1381_),
    .A2(_1417_),
    .A3(_1398_),
    .S0(net195),
    .S1(net203),
    .X(_3063_));
 sky130_fd_sc_hd__mux2_1 _5900_ (.A0(_2978_),
    .A1(_3063_),
    .S(net201),
    .X(_3064_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(_2879_),
    .A1(_3064_),
    .S(net210),
    .X(_3065_));
 sky130_fd_sc_hd__nand2_1 _5902_ (.A(_2720_),
    .B(_3065_),
    .Y(_3066_));
 sky130_fd_sc_hd__nor2_1 _5903_ (.A(net189),
    .B(_2871_),
    .Y(_3067_));
 sky130_fd_sc_hd__nor2_1 _5904_ (.A(net207),
    .B(_2865_),
    .Y(_3068_));
 sky130_fd_sc_hd__o31a_1 _5905_ (.A1(_2675_),
    .A2(_3067_),
    .A3(_3068_),
    .B1(_3066_),
    .X(_3069_));
 sky130_fd_sc_hd__o22a_1 _5906_ (.A1(net282),
    .A2(_3058_),
    .B1(_3069_),
    .B2(net212),
    .X(_3070_));
 sky130_fd_sc_hd__or3b_1 _5907_ (.A(_3061_),
    .B(_3062_),
    .C_N(_3070_),
    .X(_3071_));
 sky130_fd_sc_hd__a21o_1 _5908_ (.A1(_1354_),
    .A2(_1371_),
    .B1(net219),
    .X(_3072_));
 sky130_fd_sc_hd__and3_1 _5909_ (.A(net435),
    .B(_3071_),
    .C(_3072_),
    .X(_0637_));
 sky130_fd_sc_hd__xnor2_1 _5910_ (.A(_1387_),
    .B(net314),
    .Y(_3073_));
 sky130_fd_sc_hd__or2_1 _5911_ (.A(_1389_),
    .B(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_1389_),
    .B(_3073_),
    .Y(_3075_));
 sky130_fd_sc_hd__nand2_1 _5913_ (.A(_3074_),
    .B(_3075_),
    .Y(_3076_));
 sky130_fd_sc_hd__o21ai_2 _5914_ (.A1(_3053_),
    .A2(_3055_),
    .B1(_3056_),
    .Y(_3077_));
 sky130_fd_sc_hd__xor2_1 _5915_ (.A(_3076_),
    .B(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__a21oi_1 _5916_ (.A1(_1389_),
    .A2(net311),
    .B1(_1387_),
    .Y(_3079_));
 sky130_fd_sc_hd__o221a_1 _5917_ (.A1(_2714_),
    .A2(_3076_),
    .B1(_3079_),
    .B2(_2718_),
    .C1(_2724_),
    .X(_3080_));
 sky130_fd_sc_hd__o21a_1 _5918_ (.A1(net187),
    .A2(_2894_),
    .B1(_2986_),
    .X(_3081_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_2891_),
    .B(_2921_),
    .Y(_3082_));
 sky130_fd_sc_hd__o211a_1 _5920_ (.A1(_2672_),
    .A2(_3081_),
    .B1(_3082_),
    .C1(net211),
    .X(_3083_));
 sky130_fd_sc_hd__o21ba_1 _5921_ (.A1(net186),
    .A2(_2905_),
    .B1_N(_2675_),
    .X(_3084_));
 sky130_fd_sc_hd__o21ai_1 _5922_ (.A1(net209),
    .A2(_2889_),
    .B1(_3084_),
    .Y(_3085_));
 sky130_fd_sc_hd__mux2_1 _5923_ (.A0(_1389_),
    .A1(_1371_),
    .S(net195),
    .X(_3086_));
 sky130_fd_sc_hd__mux2_1 _5924_ (.A0(_3045_),
    .A1(_3086_),
    .S(_1449_),
    .X(_3087_));
 sky130_fd_sc_hd__inv_2 _5925_ (.A(_3087_),
    .Y(_3088_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(_2998_),
    .A1(_3087_),
    .S(net200),
    .X(_3089_));
 sky130_fd_sc_hd__nor2_1 _5927_ (.A(net188),
    .B(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__a211o_1 _5928_ (.A1(net188),
    .A2(_2902_),
    .B1(_3090_),
    .C1(_2721_),
    .X(_3091_));
 sky130_fd_sc_hd__a31o_1 _5929_ (.A1(net216),
    .A2(_3085_),
    .A3(_3091_),
    .B1(_3083_),
    .X(_3092_));
 sky130_fd_sc_hd__o211ai_1 _5930_ (.A1(_2712_),
    .A2(_3078_),
    .B1(_3080_),
    .C1(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__a21o_1 _5931_ (.A1(_1387_),
    .A2(_1389_),
    .B1(_2724_),
    .X(_3094_));
 sky130_fd_sc_hd__and3_1 _5932_ (.A(net440),
    .B(_3093_),
    .C(_3094_),
    .X(_0638_));
 sky130_fd_sc_hd__a21bo_1 _5933_ (.A1(_3074_),
    .A2(_3077_),
    .B1_N(_3075_),
    .X(_3095_));
 sky130_fd_sc_hd__xnor2_1 _5934_ (.A(_1504_),
    .B(net314),
    .Y(_3096_));
 sky130_fd_sc_hd__nor2_1 _5935_ (.A(_1506_),
    .B(_3096_),
    .Y(_3097_));
 sky130_fd_sc_hd__or2_1 _5936_ (.A(_1506_),
    .B(_3096_),
    .X(_3098_));
 sky130_fd_sc_hd__and2_1 _5937_ (.A(_1506_),
    .B(_3096_),
    .X(_3099_));
 sky130_fd_sc_hd__nor2_1 _5938_ (.A(_3097_),
    .B(_3099_),
    .Y(_3100_));
 sky130_fd_sc_hd__nor2_1 _5939_ (.A(_3095_),
    .B(_3100_),
    .Y(_3101_));
 sky130_fd_sc_hd__a21o_1 _5940_ (.A1(_3095_),
    .A2(_3100_),
    .B1(net283),
    .X(_3102_));
 sky130_fd_sc_hd__mux4_1 _5941_ (.A0(_1371_),
    .A1(_1381_),
    .A2(_1506_),
    .A3(_1389_),
    .S0(net193),
    .S1(net206),
    .X(_3103_));
 sky130_fd_sc_hd__mux2_1 _5942_ (.A0(_3024_),
    .A1(_3103_),
    .S(net200),
    .X(_3104_));
 sky130_fd_sc_hd__nor2_1 _5943_ (.A(net188),
    .B(_3104_),
    .Y(_3105_));
 sky130_fd_sc_hd__a21o_1 _5944_ (.A1(net188),
    .A2(_2933_),
    .B1(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__nor2_2 _5945_ (.A(net207),
    .B(_2919_),
    .Y(_3107_));
 sky130_fd_sc_hd__nor2_1 _5946_ (.A(net188),
    .B(_2936_),
    .Y(_3108_));
 sky130_fd_sc_hd__o32a_1 _5947_ (.A1(_2675_),
    .A2(_3107_),
    .A3(_3108_),
    .B1(_2721_),
    .B2(_3106_),
    .X(_3109_));
 sky130_fd_sc_hd__a21oi_1 _5948_ (.A1(_1506_),
    .A2(net311),
    .B1(_1504_),
    .Y(_3110_));
 sky130_fd_sc_hd__o221a_1 _5949_ (.A1(_1507_),
    .A2(_2714_),
    .B1(_2718_),
    .B2(_3110_),
    .C1(net219),
    .X(_3111_));
 sky130_fd_sc_hd__a21bo_1 _5950_ (.A1(net207),
    .A2(_2926_),
    .B1_N(_2986_),
    .X(_3112_));
 sky130_fd_sc_hd__a22o_1 _5951_ (.A1(net207),
    .A2(_2924_),
    .B1(_3112_),
    .B2(_2671_),
    .X(_3113_));
 sky130_fd_sc_hd__nand2_2 _5952_ (.A(net211),
    .B(_3113_),
    .Y(_3114_));
 sky130_fd_sc_hd__o211a_1 _5953_ (.A1(net214),
    .A2(_3109_),
    .B1(_3111_),
    .C1(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__o21ai_1 _5954_ (.A1(_3101_),
    .A2(_3102_),
    .B1(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hd__a21o_1 _5955_ (.A1(_1504_),
    .A2(_1506_),
    .B1(net219),
    .X(_3117_));
 sky130_fd_sc_hd__and3_1 _5956_ (.A(net444),
    .B(_3116_),
    .C(_3117_),
    .X(_0639_));
 sky130_fd_sc_hd__xnor2_1 _5957_ (.A(_1511_),
    .B(net314),
    .Y(_3118_));
 sky130_fd_sc_hd__nor2_1 _5958_ (.A(_1513_),
    .B(_3118_),
    .Y(_3119_));
 sky130_fd_sc_hd__nand2_1 _5959_ (.A(_1513_),
    .B(_3118_),
    .Y(_3120_));
 sky130_fd_sc_hd__nand2b_1 _5960_ (.A_N(_3119_),
    .B(_3120_),
    .Y(_3121_));
 sky130_fd_sc_hd__a21oi_1 _5961_ (.A1(_3095_),
    .A2(_3098_),
    .B1(_3099_),
    .Y(_3122_));
 sky130_fd_sc_hd__xnor2_1 _5962_ (.A(_3121_),
    .B(_3122_),
    .Y(_3123_));
 sky130_fd_sc_hd__nor2_1 _5963_ (.A(net283),
    .B(_3123_),
    .Y(_3124_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(_2955_),
    .A1(_2961_),
    .S(net186),
    .X(_3125_));
 sky130_fd_sc_hd__a21oi_4 _5965_ (.A1(net211),
    .A2(net190),
    .B1(_2672_),
    .Y(_3126_));
 sky130_fd_sc_hd__a21o_2 _5966_ (.A1(net211),
    .A2(net190),
    .B1(_2672_),
    .X(_3127_));
 sky130_fd_sc_hd__nor2_2 _5967_ (.A(net212),
    .B(_2674_),
    .Y(_3128_));
 sky130_fd_sc_hd__nor2_2 _5968_ (.A(_3126_),
    .B(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__mux2_1 _5969_ (.A0(_1513_),
    .A1(_1506_),
    .S(net195),
    .X(_3130_));
 sky130_fd_sc_hd__mux2_1 _5970_ (.A0(_3086_),
    .A1(_3130_),
    .S(net205),
    .X(_3131_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(_3046_),
    .A1(_3131_),
    .S(net200),
    .X(_3132_));
 sky130_fd_sc_hd__mux2_1 _5972_ (.A0(_2952_),
    .A1(_3132_),
    .S(net209),
    .X(_3133_));
 sky130_fd_sc_hd__a221o_1 _5973_ (.A1(_1513_),
    .A2(net311),
    .B1(net281),
    .B2(_1511_),
    .C1(net221),
    .X(_3134_));
 sky130_fd_sc_hd__nor2_1 _5974_ (.A(_2714_),
    .B(_3121_),
    .Y(_3135_));
 sky130_fd_sc_hd__and3_1 _5975_ (.A(net208),
    .B(net199),
    .C(_2830_),
    .X(_3136_));
 sky130_fd_sc_hd__a311o_1 _5976_ (.A1(net217),
    .A2(_2720_),
    .A3(_3133_),
    .B1(_3134_),
    .C1(_3135_),
    .X(_3137_));
 sky130_fd_sc_hd__o21a_1 _5977_ (.A1(net215),
    .A2(_3136_),
    .B1(_2673_),
    .X(_3138_));
 sky130_fd_sc_hd__o22a_1 _5978_ (.A1(net212),
    .A2(_3125_),
    .B1(_3126_),
    .B2(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__a21o_1 _5979_ (.A1(_1511_),
    .A2(_1513_),
    .B1(net219),
    .X(_3140_));
 sky130_fd_sc_hd__o311a_1 _5980_ (.A1(_3124_),
    .A2(_3137_),
    .A3(_3139_),
    .B1(_3140_),
    .C1(net444),
    .X(_0640_));
 sky130_fd_sc_hd__o21ai_2 _5981_ (.A1(_3119_),
    .A2(_3122_),
    .B1(_3120_),
    .Y(_3141_));
 sky130_fd_sc_hd__xnor2_1 _5982_ (.A(_1549_),
    .B(net314),
    .Y(_3142_));
 sky130_fd_sc_hd__nor2_1 _5983_ (.A(_1551_),
    .B(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__or2_1 _5984_ (.A(_1551_),
    .B(_3142_),
    .X(_3144_));
 sky130_fd_sc_hd__and2_1 _5985_ (.A(_1551_),
    .B(_3142_),
    .X(_3145_));
 sky130_fd_sc_hd__nor2_1 _5986_ (.A(_3143_),
    .B(_3145_),
    .Y(_3146_));
 sky130_fd_sc_hd__or2_1 _5987_ (.A(_3141_),
    .B(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__a21oi_1 _5988_ (.A1(_3141_),
    .A2(_3146_),
    .B1(net283),
    .Y(_3148_));
 sky130_fd_sc_hd__mux4_1 _5989_ (.A0(_1506_),
    .A1(_1551_),
    .A2(_1389_),
    .A3(_1513_),
    .S0(net206),
    .S1(net195),
    .X(_3149_));
 sky130_fd_sc_hd__mux2_1 _5990_ (.A0(_3063_),
    .A1(_3149_),
    .S(net201),
    .X(_3150_));
 sky130_fd_sc_hd__mux2_1 _5991_ (.A0(_2979_),
    .A1(_3150_),
    .S(net210),
    .X(_3151_));
 sky130_fd_sc_hd__a21oi_1 _5992_ (.A1(net214),
    .A2(_2729_),
    .B1(_2721_),
    .Y(_3152_));
 sky130_fd_sc_hd__o21a_1 _5993_ (.A1(net214),
    .A2(_3151_),
    .B1(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__o21ba_1 _5994_ (.A1(net214),
    .A2(_2705_),
    .B1_N(_3129_),
    .X(_3154_));
 sky130_fd_sc_hd__a21o_1 _5995_ (.A1(_1551_),
    .A2(_2716_),
    .B1(_1549_),
    .X(_3155_));
 sky130_fd_sc_hd__a221o_1 _5996_ (.A1(_1553_),
    .A2(_2713_),
    .B1(net281),
    .B2(_3155_),
    .C1(net221),
    .X(_3156_));
 sky130_fd_sc_hd__or3_1 _5997_ (.A(_3153_),
    .B(_3154_),
    .C(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__a21o_1 _5998_ (.A1(_3147_),
    .A2(_3148_),
    .B1(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__a21o_1 _5999_ (.A1(_1549_),
    .A2(net2258),
    .B1(_2724_),
    .X(_3159_));
 sky130_fd_sc_hd__and3_1 _6000_ (.A(net444),
    .B(_3158_),
    .C(net2259),
    .X(_0641_));
 sky130_fd_sc_hd__xnor2_1 _6001_ (.A(_1557_),
    .B(_2708_),
    .Y(_3160_));
 sky130_fd_sc_hd__or2_1 _6002_ (.A(_1559_),
    .B(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__nand2_1 _6003_ (.A(_1559_),
    .B(_3160_),
    .Y(_3162_));
 sky130_fd_sc_hd__nand2_1 _6004_ (.A(_3161_),
    .B(_3162_),
    .Y(_3163_));
 sky130_fd_sc_hd__a21o_1 _6005_ (.A1(_3141_),
    .A2(_3144_),
    .B1(_3145_),
    .X(_3164_));
 sky130_fd_sc_hd__xor2_1 _6006_ (.A(_3163_),
    .B(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__or2_1 _6007_ (.A(net205),
    .B(_3130_),
    .X(_3166_));
 sky130_fd_sc_hd__mux2_1 _6008_ (.A0(_1559_),
    .A1(_1551_),
    .S(net193),
    .X(_3167_));
 sky130_fd_sc_hd__o21ai_1 _6009_ (.A1(net202),
    .A2(_3167_),
    .B1(_3166_),
    .Y(_3168_));
 sky130_fd_sc_hd__mux2_1 _6010_ (.A0(_3088_),
    .A1(_3168_),
    .S(net200),
    .X(_3169_));
 sky130_fd_sc_hd__nand2_1 _6011_ (.A(net189),
    .B(_2999_),
    .Y(_3170_));
 sky130_fd_sc_hd__o211a_1 _6012_ (.A1(net189),
    .A2(_3169_),
    .B1(_3170_),
    .C1(net216),
    .X(_3171_));
 sky130_fd_sc_hd__a211o_1 _6013_ (.A1(net214),
    .A2(_2763_),
    .B1(_3171_),
    .C1(_2721_),
    .X(_3172_));
 sky130_fd_sc_hd__o2bb2a_1 _6014_ (.A1_N(_1559_),
    .A2_N(_2716_),
    .B1(_2718_),
    .B2(_1557_),
    .X(_3173_));
 sky130_fd_sc_hd__o2bb2a_1 _6015_ (.A1_N(_2747_),
    .A2_N(_3128_),
    .B1(_3163_),
    .B2(net312),
    .X(_3174_));
 sky130_fd_sc_hd__and3_1 _6016_ (.A(_2724_),
    .B(_3173_),
    .C(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__nor2_1 _6017_ (.A(net212),
    .B(_2744_),
    .Y(_3176_));
 sky130_fd_sc_hd__o221a_1 _6018_ (.A1(net283),
    .A2(_3165_),
    .B1(_3176_),
    .B2(_3127_),
    .C1(_3175_),
    .X(_3177_));
 sky130_fd_sc_hd__nand2b_1 _6019_ (.A_N(_1557_),
    .B(_1559_),
    .Y(_3178_));
 sky130_fd_sc_hd__a221oi_1 _6020_ (.A1(_3172_),
    .A2(_3177_),
    .B1(_3178_),
    .B2(net220),
    .C1(net63),
    .Y(_0642_));
 sky130_fd_sc_hd__a21bo_1 _6021_ (.A1(_3161_),
    .A2(_3164_),
    .B1_N(_3162_),
    .X(_3179_));
 sky130_fd_sc_hd__xnor2_1 _6022_ (.A(_1582_),
    .B(net314),
    .Y(_3180_));
 sky130_fd_sc_hd__nor2_1 _6023_ (.A(_1584_),
    .B(_3180_),
    .Y(_3181_));
 sky130_fd_sc_hd__or2_1 _6024_ (.A(_1584_),
    .B(_3180_),
    .X(_3182_));
 sky130_fd_sc_hd__and2_1 _6025_ (.A(_1584_),
    .B(_3180_),
    .X(_3183_));
 sky130_fd_sc_hd__nor2_1 _6026_ (.A(_3181_),
    .B(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__xnor2_1 _6027_ (.A(_3179_),
    .B(_3184_),
    .Y(_3185_));
 sky130_fd_sc_hd__a2111oi_1 _6028_ (.A1(net212),
    .A2(net190),
    .B1(_2672_),
    .C1(_2806_),
    .D1(_2812_),
    .Y(_3186_));
 sky130_fd_sc_hd__nand2_2 _6029_ (.A(_1638_),
    .B(_2671_),
    .Y(_3187_));
 sky130_fd_sc_hd__a21oi_1 _6030_ (.A1(_2791_),
    .A2(_3187_),
    .B1(net217),
    .Y(_3188_));
 sky130_fd_sc_hd__a221o_1 _6031_ (.A1(_1584_),
    .A2(net311),
    .B1(net281),
    .B2(_1582_),
    .C1(net221),
    .X(_3189_));
 sky130_fd_sc_hd__a2111o_1 _6032_ (.A1(_1585_),
    .A2(_2713_),
    .B1(net185),
    .C1(_3188_),
    .D1(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__mux4_1 _6033_ (.A0(_1551_),
    .A1(_1584_),
    .A2(_1513_),
    .A3(_1559_),
    .S0(net205),
    .S1(net193),
    .X(_3191_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(_3103_),
    .A1(_3191_),
    .S(net200),
    .X(_3192_));
 sky130_fd_sc_hd__mux2_1 _6035_ (.A0(_3025_),
    .A1(_3192_),
    .S(net209),
    .X(_3193_));
 sky130_fd_sc_hd__a21bo_1 _6036_ (.A1(_2720_),
    .A2(_3193_),
    .B1_N(_2815_),
    .X(_3194_));
 sky130_fd_sc_hd__a2bb2o_1 _6037_ (.A1_N(_2712_),
    .A2_N(_3185_),
    .B1(_3194_),
    .B2(net216),
    .X(_3195_));
 sky130_fd_sc_hd__a21o_1 _6038_ (.A1(_1582_),
    .A2(_1584_),
    .B1(_2724_),
    .X(_3196_));
 sky130_fd_sc_hd__o211a_1 _6039_ (.A1(_3190_),
    .A2(_3195_),
    .B1(_3196_),
    .C1(net438),
    .X(_0643_));
 sky130_fd_sc_hd__xnor2_1 _6040_ (.A(_1564_),
    .B(_2708_),
    .Y(_3197_));
 sky130_fd_sc_hd__or2_1 _6041_ (.A(_1566_),
    .B(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_1566_),
    .B(_3197_),
    .Y(_3199_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_3198_),
    .B(_3199_),
    .Y(_3200_));
 sky130_fd_sc_hd__a21o_1 _6044_ (.A1(_3179_),
    .A2(_3182_),
    .B1(_3183_),
    .X(_3201_));
 sky130_fd_sc_hd__xor2_1 _6045_ (.A(_3200_),
    .B(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__mux2_1 _6046_ (.A0(_1566_),
    .A1(_1584_),
    .S(net193),
    .X(_3203_));
 sky130_fd_sc_hd__mux2_1 _6047_ (.A0(_3167_),
    .A1(_3203_),
    .S(net205),
    .X(_3204_));
 sky130_fd_sc_hd__mux2_1 _6048_ (.A0(_3131_),
    .A1(_3204_),
    .S(net200),
    .X(_3205_));
 sky130_fd_sc_hd__mux2_1 _6049_ (.A0(_3047_),
    .A1(_3205_),
    .S(net209),
    .X(_3206_));
 sky130_fd_sc_hd__a31o_1 _6050_ (.A1(net209),
    .A2(net200),
    .A3(_2842_),
    .B1(net215),
    .X(_3207_));
 sky130_fd_sc_hd__o211a_1 _6051_ (.A1(net212),
    .A2(_3206_),
    .B1(_3207_),
    .C1(_2720_),
    .X(_3208_));
 sky130_fd_sc_hd__nand2_1 _6052_ (.A(_2832_),
    .B(_3128_),
    .Y(_3209_));
 sky130_fd_sc_hd__a21oi_1 _6053_ (.A1(_1566_),
    .A2(net310),
    .B1(net220),
    .Y(_3210_));
 sky130_fd_sc_hd__o221a_1 _6054_ (.A1(_1564_),
    .A2(_2718_),
    .B1(_3200_),
    .B2(net312),
    .C1(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__o21ai_1 _6055_ (.A1(net212),
    .A2(_2829_),
    .B1(_3126_),
    .Y(_3212_));
 sky130_fd_sc_hd__and4b_1 _6056_ (.A_N(_3208_),
    .B(_3209_),
    .C(_3211_),
    .D(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__o21ai_1 _6057_ (.A1(net282),
    .A2(_3202_),
    .B1(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__and2b_1 _6058_ (.A_N(_1564_),
    .B(_1566_),
    .X(_3215_));
 sky130_fd_sc_hd__o211a_1 _6059_ (.A1(net219),
    .A2(_3215_),
    .B1(_3214_),
    .C1(net438),
    .X(_0644_));
 sky130_fd_sc_hd__a21bo_1 _6060_ (.A1(_3198_),
    .A2(_3201_),
    .B1_N(_3199_),
    .X(_3216_));
 sky130_fd_sc_hd__xnor2_1 _6061_ (.A(_1573_),
    .B(net313),
    .Y(_3217_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(_1575_),
    .B(_3217_),
    .Y(_3218_));
 sky130_fd_sc_hd__or2_1 _6063_ (.A(_1575_),
    .B(_3217_),
    .X(_3219_));
 sky130_fd_sc_hd__and2_1 _6064_ (.A(_1575_),
    .B(_3217_),
    .X(_3220_));
 sky130_fd_sc_hd__nor2_1 _6065_ (.A(_3218_),
    .B(_3220_),
    .Y(_3221_));
 sky130_fd_sc_hd__a21oi_1 _6066_ (.A1(_3216_),
    .A2(_3221_),
    .B1(net283),
    .Y(_3222_));
 sky130_fd_sc_hd__o21a_1 _6067_ (.A1(_3216_),
    .A2(_3221_),
    .B1(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__mux4_1 _6068_ (.A0(_1575_),
    .A1(_1584_),
    .A2(_1566_),
    .A3(_1559_),
    .S0(net203),
    .S1(net195),
    .X(_3224_));
 sky130_fd_sc_hd__mux2_1 _6069_ (.A0(_3149_),
    .A1(_3224_),
    .S(net201),
    .X(_3225_));
 sky130_fd_sc_hd__mux2_1 _6070_ (.A0(_3064_),
    .A1(_3225_),
    .S(net210),
    .X(_3226_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(net214),
    .B(_2880_),
    .Y(_3227_));
 sky130_fd_sc_hd__o211a_1 _6072_ (.A1(net214),
    .A2(_3226_),
    .B1(_3227_),
    .C1(_2720_),
    .X(_3228_));
 sky130_fd_sc_hd__a21o_1 _6073_ (.A1(_1575_),
    .A2(net311),
    .B1(_1573_),
    .X(_3229_));
 sky130_fd_sc_hd__a221o_1 _6074_ (.A1(_1577_),
    .A2(_2713_),
    .B1(net281),
    .B2(_3229_),
    .C1(net220),
    .X(_3230_));
 sky130_fd_sc_hd__o21a_1 _6075_ (.A1(net208),
    .A2(_2867_),
    .B1(_3128_),
    .X(_3231_));
 sky130_fd_sc_hd__o22a_1 _6076_ (.A1(net212),
    .A2(_2869_),
    .B1(_3126_),
    .B2(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__or4_1 _6077_ (.A(_3223_),
    .B(_3228_),
    .C(_3230_),
    .D(_3232_),
    .X(_3233_));
 sky130_fd_sc_hd__a21o_1 _6078_ (.A1(_1573_),
    .A2(_1575_),
    .B1(net219),
    .X(_3234_));
 sky130_fd_sc_hd__and3_1 _6079_ (.A(net436),
    .B(_3233_),
    .C(_3234_),
    .X(_0645_));
 sky130_fd_sc_hd__xnor2_1 _6080_ (.A(_1539_),
    .B(net313),
    .Y(_3235_));
 sky130_fd_sc_hd__or2_1 _6081_ (.A(_1541_),
    .B(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__nand2_1 _6082_ (.A(_1541_),
    .B(_3235_),
    .Y(_3237_));
 sky130_fd_sc_hd__nand2_1 _6083_ (.A(_3236_),
    .B(_3237_),
    .Y(_3238_));
 sky130_fd_sc_hd__a21o_1 _6084_ (.A1(_3216_),
    .A2(_3219_),
    .B1(_3220_),
    .X(_3239_));
 sky130_fd_sc_hd__nand2_1 _6085_ (.A(_3238_),
    .B(_3239_),
    .Y(_3240_));
 sky130_fd_sc_hd__or2_1 _6086_ (.A(_3238_),
    .B(_3239_),
    .X(_3241_));
 sky130_fd_sc_hd__a21oi_1 _6087_ (.A1(_3240_),
    .A2(_3241_),
    .B1(net282),
    .Y(_3242_));
 sky130_fd_sc_hd__o21a_1 _6088_ (.A1(net211),
    .A2(_2895_),
    .B1(_3126_),
    .X(_3243_));
 sky130_fd_sc_hd__a221o_1 _6089_ (.A1(_1541_),
    .A2(net310),
    .B1(net281),
    .B2(_1539_),
    .C1(net220),
    .X(_3244_));
 sky130_fd_sc_hd__o22a_1 _6090_ (.A1(net211),
    .A2(_2893_),
    .B1(_3238_),
    .B2(net312),
    .X(_3245_));
 sky130_fd_sc_hd__nand2_1 _6091_ (.A(net186),
    .B(_3089_),
    .Y(_3246_));
 sky130_fd_sc_hd__mux2_1 _6092_ (.A0(_1541_),
    .A1(_1575_),
    .S(net192),
    .X(_3247_));
 sky130_fd_sc_hd__mux2_1 _6093_ (.A0(_3203_),
    .A1(_3247_),
    .S(net206),
    .X(_3248_));
 sky130_fd_sc_hd__inv_2 _6094_ (.A(_3248_),
    .Y(_3249_));
 sky130_fd_sc_hd__mux2_1 _6095_ (.A0(_3168_),
    .A1(_3249_),
    .S(net199),
    .X(_3250_));
 sky130_fd_sc_hd__o211a_1 _6096_ (.A1(net186),
    .A2(_3250_),
    .B1(_3246_),
    .C1(net216),
    .X(_3251_));
 sky130_fd_sc_hd__a21oi_1 _6097_ (.A1(_2727_),
    .A2(_2903_),
    .B1(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hd__or4b_1 _6098_ (.A(_3243_),
    .B(_3244_),
    .C(_3252_),
    .D_N(_3245_),
    .X(_3253_));
 sky130_fd_sc_hd__a21o_1 _6099_ (.A1(_1539_),
    .A2(_1541_),
    .B1(net218),
    .X(_3254_));
 sky130_fd_sc_hd__o211a_1 _6100_ (.A1(_3242_),
    .A2(_3253_),
    .B1(_3254_),
    .C1(net436),
    .X(_0646_));
 sky130_fd_sc_hd__a21bo_1 _6101_ (.A1(_3236_),
    .A2(_3239_),
    .B1_N(_3237_),
    .X(_3255_));
 sky130_fd_sc_hd__xnor2_1 _6102_ (.A(_1522_),
    .B(net313),
    .Y(_3256_));
 sky130_fd_sc_hd__nor2_1 _6103_ (.A(_1524_),
    .B(_3256_),
    .Y(_3257_));
 sky130_fd_sc_hd__or2_1 _6104_ (.A(_1524_),
    .B(_3256_),
    .X(_3258_));
 sky130_fd_sc_hd__and2_1 _6105_ (.A(_1524_),
    .B(_3256_),
    .X(_3259_));
 sky130_fd_sc_hd__nor2_1 _6106_ (.A(_3257_),
    .B(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__xnor2_1 _6107_ (.A(_3255_),
    .B(_3260_),
    .Y(_3261_));
 sky130_fd_sc_hd__o211a_1 _6108_ (.A1(net207),
    .A2(_2926_),
    .B1(_3126_),
    .C1(_2920_),
    .X(_3262_));
 sky130_fd_sc_hd__a21o_1 _6109_ (.A1(_1524_),
    .A2(net310),
    .B1(_1522_),
    .X(_3263_));
 sky130_fd_sc_hd__a221o_1 _6110_ (.A1(_1525_),
    .A2(_2713_),
    .B1(net281),
    .B2(_3263_),
    .C1(net220),
    .X(_3264_));
 sky130_fd_sc_hd__a21oi_1 _6111_ (.A1(_2934_),
    .A2(_3187_),
    .B1(net215),
    .Y(_3265_));
 sky130_fd_sc_hd__mux4_1 _6112_ (.A0(_1524_),
    .A1(_1541_),
    .A2(_1575_),
    .A3(_1566_),
    .S0(net192),
    .S1(net202),
    .X(_3266_));
 sky130_fd_sc_hd__mux2_1 _6113_ (.A0(_3191_),
    .A1(_3266_),
    .S(net199),
    .X(_3267_));
 sky130_fd_sc_hd__mux2_1 _6114_ (.A0(_3104_),
    .A1(_3267_),
    .S(net207),
    .X(_3268_));
 sky130_fd_sc_hd__a21o_1 _6115_ (.A1(_2720_),
    .A2(_3268_),
    .B1(_2925_),
    .X(_3269_));
 sky130_fd_sc_hd__a2bb2o_1 _6116_ (.A1_N(net282),
    .A2_N(_3261_),
    .B1(_3269_),
    .B2(net215),
    .X(_3270_));
 sky130_fd_sc_hd__or4_1 _6117_ (.A(_3262_),
    .B(_3264_),
    .C(_3265_),
    .D(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__a21o_1 _6118_ (.A1(_1522_),
    .A2(net2324),
    .B1(net219),
    .X(_3272_));
 sky130_fd_sc_hd__and3_1 _6119_ (.A(net436),
    .B(_3271_),
    .C(_3272_),
    .X(_0647_));
 sky130_fd_sc_hd__xnor2_1 _6120_ (.A(_1530_),
    .B(net316),
    .Y(_3273_));
 sky130_fd_sc_hd__or2_1 _6121_ (.A(_1533_),
    .B(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__and2_1 _6122_ (.A(_1533_),
    .B(_3273_),
    .X(_3275_));
 sky130_fd_sc_hd__nand2_1 _6123_ (.A(_1533_),
    .B(_3273_),
    .Y(_3276_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(_3274_),
    .B(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__a21o_1 _6125_ (.A1(_3255_),
    .A2(_3258_),
    .B1(_3259_),
    .X(_3278_));
 sky130_fd_sc_hd__xor2_1 _6126_ (.A(_3277_),
    .B(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__a21oi_1 _6127_ (.A1(_1533_),
    .A2(net310),
    .B1(_1531_),
    .Y(_3280_));
 sky130_fd_sc_hd__o221ai_2 _6128_ (.A1(net312),
    .A2(_3277_),
    .B1(_3280_),
    .B2(_2718_),
    .C1(net218),
    .Y(_3281_));
 sky130_fd_sc_hd__a21oi_1 _6129_ (.A1(_2953_),
    .A2(_3187_),
    .B1(net215),
    .Y(_3282_));
 sky130_fd_sc_hd__a211o_1 _6130_ (.A1(_2965_),
    .A2(_3126_),
    .B1(_3281_),
    .C1(_3282_),
    .X(_3283_));
 sky130_fd_sc_hd__mux2_1 _6131_ (.A0(_1533_),
    .A1(_1524_),
    .S(net191),
    .X(_3284_));
 sky130_fd_sc_hd__mux2_1 _6132_ (.A0(_3247_),
    .A1(_3284_),
    .S(net205),
    .X(_3285_));
 sky130_fd_sc_hd__mux2_1 _6133_ (.A0(_3204_),
    .A1(_3285_),
    .S(net199),
    .X(_3286_));
 sky130_fd_sc_hd__mux2_1 _6134_ (.A0(_3132_),
    .A1(_3286_),
    .S(net207),
    .X(_3287_));
 sky130_fd_sc_hd__a21o_1 _6135_ (.A1(_2720_),
    .A2(_3287_),
    .B1(_2964_),
    .X(_3288_));
 sky130_fd_sc_hd__a2bb2o_1 _6136_ (.A1_N(net282),
    .A2_N(_3279_),
    .B1(_3288_),
    .B2(net215),
    .X(_3289_));
 sky130_fd_sc_hd__a21o_1 _6137_ (.A1(_1531_),
    .A2(_1533_),
    .B1(net218),
    .X(_3290_));
 sky130_fd_sc_hd__o211a_1 _6138_ (.A1(_3283_),
    .A2(_3289_),
    .B1(_3290_),
    .C1(net435),
    .X(_0648_));
 sky130_fd_sc_hd__a21o_1 _6139_ (.A1(_3274_),
    .A2(_3278_),
    .B1(_3275_),
    .X(_3291_));
 sky130_fd_sc_hd__xnor2_1 _6140_ (.A(_1646_),
    .B(net313),
    .Y(_3292_));
 sky130_fd_sc_hd__nor2_1 _6141_ (.A(_1648_),
    .B(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__or2_1 _6142_ (.A(_1648_),
    .B(_3292_),
    .X(_3294_));
 sky130_fd_sc_hd__and2_1 _6143_ (.A(_1648_),
    .B(_3292_),
    .X(_3295_));
 sky130_fd_sc_hd__nor2_1 _6144_ (.A(_3293_),
    .B(_3295_),
    .Y(_3296_));
 sky130_fd_sc_hd__nor2_1 _6145_ (.A(_3291_),
    .B(_3296_),
    .Y(_3297_));
 sky130_fd_sc_hd__a21o_1 _6146_ (.A1(_3291_),
    .A2(_3296_),
    .B1(net282),
    .X(_3298_));
 sky130_fd_sc_hd__mux4_2 _6147_ (.A0(_1524_),
    .A1(_1541_),
    .A2(_1648_),
    .A3(_1533_),
    .S0(net192),
    .S1(net205),
    .X(_3299_));
 sky130_fd_sc_hd__mux2_1 _6148_ (.A0(_3224_),
    .A1(_3299_),
    .S(net201),
    .X(_3300_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(_3150_),
    .A1(_3300_),
    .S(net210),
    .X(_3301_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(net214),
    .B(_2981_),
    .Y(_3302_));
 sky130_fd_sc_hd__o211a_1 _6151_ (.A1(net214),
    .A2(_3301_),
    .B1(_3302_),
    .C1(_2720_),
    .X(_3303_));
 sky130_fd_sc_hd__a221o_1 _6152_ (.A1(_1648_),
    .A2(net310),
    .B1(net281),
    .B2(_1646_),
    .C1(net220),
    .X(_3304_));
 sky130_fd_sc_hd__a21oi_1 _6153_ (.A1(net215),
    .A2(_2986_),
    .B1(_3127_),
    .Y(_3305_));
 sky130_fd_sc_hd__nor2_1 _6154_ (.A(_3304_),
    .B(_3305_),
    .Y(_3306_));
 sky130_fd_sc_hd__o221a_1 _6155_ (.A1(_1650_),
    .A2(net312),
    .B1(_2985_),
    .B2(_3129_),
    .C1(_3306_),
    .X(_3307_));
 sky130_fd_sc_hd__o21ai_1 _6156_ (.A1(_3297_),
    .A2(_3298_),
    .B1(_3307_),
    .Y(_3308_));
 sky130_fd_sc_hd__a21o_1 _6157_ (.A1(_1646_),
    .A2(net2331),
    .B1(net219),
    .X(_3309_));
 sky130_fd_sc_hd__o211a_1 _6158_ (.A1(_3303_),
    .A2(_3308_),
    .B1(net2332),
    .C1(net435),
    .X(_0649_));
 sky130_fd_sc_hd__xnor2_1 _6159_ (.A(_1616_),
    .B(net316),
    .Y(_3310_));
 sky130_fd_sc_hd__nor2_1 _6160_ (.A(_1618_),
    .B(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hd__nand2_1 _6161_ (.A(_1618_),
    .B(_3310_),
    .Y(_3312_));
 sky130_fd_sc_hd__nand2b_1 _6162_ (.A_N(_3311_),
    .B(_3312_),
    .Y(_3313_));
 sky130_fd_sc_hd__a21oi_2 _6163_ (.A1(_3291_),
    .A2(_3294_),
    .B1(_3295_),
    .Y(_3314_));
 sky130_fd_sc_hd__nor2_1 _6164_ (.A(_3313_),
    .B(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__a21o_1 _6165_ (.A1(_3313_),
    .A2(_3314_),
    .B1(net282),
    .X(_3316_));
 sky130_fd_sc_hd__nor2_1 _6166_ (.A(net209),
    .B(_3169_),
    .Y(_3317_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(_1618_),
    .A1(_1648_),
    .S(net192),
    .X(_3318_));
 sky130_fd_sc_hd__mux2_1 _6168_ (.A0(_3284_),
    .A1(_3318_),
    .S(net205),
    .X(_3319_));
 sky130_fd_sc_hd__mux2_1 _6169_ (.A0(_3248_),
    .A1(_3319_),
    .S(net199),
    .X(_3320_));
 sky130_fd_sc_hd__a211o_1 _6170_ (.A1(net209),
    .A2(_3320_),
    .B1(_3317_),
    .C1(net213),
    .X(_3321_));
 sky130_fd_sc_hd__o211a_1 _6171_ (.A1(net216),
    .A2(_3000_),
    .B1(_3321_),
    .C1(_2720_),
    .X(_3322_));
 sky130_fd_sc_hd__a21o_1 _6172_ (.A1(net215),
    .A2(_3006_),
    .B1(_3127_),
    .X(_3323_));
 sky130_fd_sc_hd__a21boi_1 _6173_ (.A1(_1618_),
    .A2(net310),
    .B1_N(_1616_),
    .Y(_3324_));
 sky130_fd_sc_hd__o221a_1 _6174_ (.A1(net312),
    .A2(_3313_),
    .B1(_3324_),
    .B2(_2718_),
    .C1(net218),
    .X(_3325_));
 sky130_fd_sc_hd__o311a_1 _6175_ (.A1(net211),
    .A2(_2746_),
    .A3(_2922_),
    .B1(_3323_),
    .C1(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__o21ai_1 _6176_ (.A1(_3315_),
    .A2(_3316_),
    .B1(_3326_),
    .Y(_3327_));
 sky130_fd_sc_hd__and2b_1 _6177_ (.A_N(_1616_),
    .B(_1618_),
    .X(_3328_));
 sky130_fd_sc_hd__o221a_1 _6178_ (.A1(_3322_),
    .A2(_3327_),
    .B1(_3328_),
    .B2(net218),
    .C1(net435),
    .X(_0650_));
 sky130_fd_sc_hd__o21ai_2 _6179_ (.A1(_3311_),
    .A2(_3314_),
    .B1(_3312_),
    .Y(_3329_));
 sky130_fd_sc_hd__xnor2_1 _6180_ (.A(_1608_),
    .B(net313),
    .Y(_3330_));
 sky130_fd_sc_hd__nor2_1 _6181_ (.A(_1611_),
    .B(_3330_),
    .Y(_3331_));
 sky130_fd_sc_hd__or2_1 _6182_ (.A(_1611_),
    .B(_3330_),
    .X(_3332_));
 sky130_fd_sc_hd__and2_1 _6183_ (.A(_1611_),
    .B(_3330_),
    .X(_3333_));
 sky130_fd_sc_hd__nor2_1 _6184_ (.A(_3331_),
    .B(_3333_),
    .Y(_3334_));
 sky130_fd_sc_hd__a21oi_1 _6185_ (.A1(_3329_),
    .A2(_3334_),
    .B1(net282),
    .Y(_3335_));
 sky130_fd_sc_hd__o21a_1 _6186_ (.A1(_3329_),
    .A2(_3334_),
    .B1(_3335_),
    .X(_3336_));
 sky130_fd_sc_hd__mux4_1 _6187_ (.A0(_1611_),
    .A1(_1618_),
    .A2(_1648_),
    .A3(_1533_),
    .S0(net191),
    .S1(net202),
    .X(_3337_));
 sky130_fd_sc_hd__mux2_1 _6188_ (.A0(_3266_),
    .A1(_3337_),
    .S(net199),
    .X(_3338_));
 sky130_fd_sc_hd__mux2_1 _6189_ (.A0(_3192_),
    .A1(_3338_),
    .S(net209),
    .X(_3339_));
 sky130_fd_sc_hd__o2bb2a_1 _6190_ (.A1_N(_2727_),
    .A2_N(_3027_),
    .B1(_3339_),
    .B2(net212),
    .X(_3340_));
 sky130_fd_sc_hd__a21oi_1 _6191_ (.A1(net215),
    .A2(_3019_),
    .B1(_3127_),
    .Y(_3341_));
 sky130_fd_sc_hd__a21o_1 _6192_ (.A1(_1611_),
    .A2(net310),
    .B1(_1608_),
    .X(_3342_));
 sky130_fd_sc_hd__a221o_1 _6193_ (.A1(_1612_),
    .A2(_2713_),
    .B1(net281),
    .B2(_3342_),
    .C1(net220),
    .X(_3343_));
 sky130_fd_sc_hd__nor2_1 _6194_ (.A(net213),
    .B(_3018_),
    .Y(_3344_));
 sky130_fd_sc_hd__or4_1 _6195_ (.A(_3340_),
    .B(_3341_),
    .C(_3343_),
    .D(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__a21o_1 _6196_ (.A1(_1608_),
    .A2(net2321),
    .B1(net218),
    .X(_3346_));
 sky130_fd_sc_hd__o211a_1 _6197_ (.A1(_3336_),
    .A2(_3345_),
    .B1(_3346_),
    .C1(net429),
    .X(_0651_));
 sky130_fd_sc_hd__xnor2_1 _6198_ (.A(_1625_),
    .B(net313),
    .Y(_3347_));
 sky130_fd_sc_hd__or2_1 _6199_ (.A(_1627_),
    .B(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__and2_1 _6200_ (.A(_1627_),
    .B(_3347_),
    .X(_3349_));
 sky130_fd_sc_hd__inv_2 _6201_ (.A(_3349_),
    .Y(_3350_));
 sky130_fd_sc_hd__nand2_1 _6202_ (.A(_3348_),
    .B(_3350_),
    .Y(_3351_));
 sky130_fd_sc_hd__a21o_1 _6203_ (.A1(_3329_),
    .A2(_3332_),
    .B1(_3333_),
    .X(_3352_));
 sky130_fd_sc_hd__xor2_1 _6204_ (.A(_3351_),
    .B(_3352_),
    .X(_3353_));
 sky130_fd_sc_hd__mux2_1 _6205_ (.A0(_1627_),
    .A1(_1611_),
    .S(net192),
    .X(_3354_));
 sky130_fd_sc_hd__mux2_1 _6206_ (.A0(_3318_),
    .A1(_3354_),
    .S(net205),
    .X(_3355_));
 sky130_fd_sc_hd__mux2_1 _6207_ (.A0(_3285_),
    .A1(_3355_),
    .S(net199),
    .X(_3356_));
 sky130_fd_sc_hd__mux2_1 _6208_ (.A0(_3205_),
    .A1(_3356_),
    .S(net210),
    .X(_3357_));
 sky130_fd_sc_hd__o2bb2a_1 _6209_ (.A1_N(_2727_),
    .A2_N(_3049_),
    .B1(_3357_),
    .B2(net212),
    .X(_3358_));
 sky130_fd_sc_hd__a21o_1 _6210_ (.A1(net215),
    .A2(_3041_),
    .B1(_3127_),
    .X(_3359_));
 sky130_fd_sc_hd__a21oi_1 _6211_ (.A1(_1627_),
    .A2(net310),
    .B1(_1625_),
    .Y(_3360_));
 sky130_fd_sc_hd__o221a_1 _6212_ (.A1(net312),
    .A2(_3351_),
    .B1(_3360_),
    .B2(_2718_),
    .C1(net218),
    .X(_3361_));
 sky130_fd_sc_hd__o311a_1 _6213_ (.A1(net211),
    .A2(_2831_),
    .A3(_2922_),
    .B1(_3359_),
    .C1(_3361_),
    .X(_3362_));
 sky130_fd_sc_hd__o21ai_1 _6214_ (.A1(net282),
    .A2(_3353_),
    .B1(_3362_),
    .Y(_3363_));
 sky130_fd_sc_hd__a21o_1 _6215_ (.A1(_1625_),
    .A2(_1627_),
    .B1(net218),
    .X(_3364_));
 sky130_fd_sc_hd__o211a_1 _6216_ (.A1(_3358_),
    .A2(_3363_),
    .B1(_3364_),
    .C1(net435),
    .X(_0652_));
 sky130_fd_sc_hd__a21oi_2 _6217_ (.A1(_3348_),
    .A2(_3352_),
    .B1(_3349_),
    .Y(_3365_));
 sky130_fd_sc_hd__xnor2_1 _6218_ (.A(_1654_),
    .B(net313),
    .Y(_3366_));
 sky130_fd_sc_hd__nor2_1 _6219_ (.A(_1656_),
    .B(_3366_),
    .Y(_3367_));
 sky130_fd_sc_hd__nand2_1 _6220_ (.A(_1656_),
    .B(_3366_),
    .Y(_3368_));
 sky130_fd_sc_hd__and2b_1 _6221_ (.A_N(_3367_),
    .B(_3368_),
    .X(_3369_));
 sky130_fd_sc_hd__xnor2_1 _6222_ (.A(_3365_),
    .B(_3369_),
    .Y(_3370_));
 sky130_fd_sc_hd__and2b_1 _6223_ (.A_N(net282),
    .B(_3370_),
    .X(_3371_));
 sky130_fd_sc_hd__mux4_1 _6224_ (.A0(_1611_),
    .A1(_1618_),
    .A2(_1656_),
    .A3(_1627_),
    .S0(net191),
    .S1(net205),
    .X(_3372_));
 sky130_fd_sc_hd__mux2_1 _6225_ (.A0(_3299_),
    .A1(_3372_),
    .S(net199),
    .X(_3373_));
 sky130_fd_sc_hd__mux2_1 _6226_ (.A0(_3225_),
    .A1(_3373_),
    .S(net209),
    .X(_3374_));
 sky130_fd_sc_hd__o2bb2a_1 _6227_ (.A1_N(_2727_),
    .A2_N(_3066_),
    .B1(_3374_),
    .B2(net213),
    .X(_3375_));
 sky130_fd_sc_hd__a21oi_1 _6228_ (.A1(net215),
    .A2(_3059_),
    .B1(_3127_),
    .Y(_3376_));
 sky130_fd_sc_hd__and3_1 _6229_ (.A(net215),
    .B(_2867_),
    .C(_2921_),
    .X(_3377_));
 sky130_fd_sc_hd__a221o_1 _6230_ (.A1(_1656_),
    .A2(net310),
    .B1(net281),
    .B2(_1654_),
    .C1(net220),
    .X(_3378_));
 sky130_fd_sc_hd__a2111o_1 _6231_ (.A1(_1658_),
    .A2(_2713_),
    .B1(_3376_),
    .C1(_3377_),
    .D1(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__a21o_1 _6232_ (.A1(_1654_),
    .A2(_1656_),
    .B1(net218),
    .X(_3380_));
 sky130_fd_sc_hd__o311a_1 _6233_ (.A1(_3371_),
    .A2(_3375_),
    .A3(_3379_),
    .B1(_3380_),
    .C1(net435),
    .X(_0653_));
 sky130_fd_sc_hd__xnor2_1 _6234_ (.A(_1600_),
    .B(net316),
    .Y(_3381_));
 sky130_fd_sc_hd__or2_1 _6235_ (.A(_1603_),
    .B(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__nand2_1 _6236_ (.A(_1603_),
    .B(_3381_),
    .Y(_3383_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_3382_),
    .B(_3383_),
    .Y(_3384_));
 sky130_fd_sc_hd__o21ai_2 _6238_ (.A1(_3365_),
    .A2(_3367_),
    .B1(_3368_),
    .Y(_3385_));
 sky130_fd_sc_hd__xor2_1 _6239_ (.A(_3384_),
    .B(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__a21o_1 _6240_ (.A1(net191),
    .A2(_1656_),
    .B1(_2739_),
    .X(_3387_));
 sky130_fd_sc_hd__mux2_1 _6241_ (.A0(_3354_),
    .A1(_3387_),
    .S(net205),
    .X(_3388_));
 sky130_fd_sc_hd__nand2_1 _6242_ (.A(net197),
    .B(_3319_),
    .Y(_3389_));
 sky130_fd_sc_hd__a21oi_1 _6243_ (.A1(net199),
    .A2(_3388_),
    .B1(net186),
    .Y(_3390_));
 sky130_fd_sc_hd__a22o_1 _6244_ (.A1(net186),
    .A2(_3250_),
    .B1(_3389_),
    .B2(_3390_),
    .X(_3391_));
 sky130_fd_sc_hd__a22o_1 _6245_ (.A1(_2727_),
    .A2(_3091_),
    .B1(_3391_),
    .B2(net216),
    .X(_3392_));
 sky130_fd_sc_hd__a21o_1 _6246_ (.A1(net215),
    .A2(_3081_),
    .B1(_3127_),
    .X(_3393_));
 sky130_fd_sc_hd__a21oi_1 _6247_ (.A1(_1603_),
    .A2(net310),
    .B1(_1601_),
    .Y(_3394_));
 sky130_fd_sc_hd__o221a_1 _6248_ (.A1(net312),
    .A2(_3384_),
    .B1(_3394_),
    .B2(_2718_),
    .C1(net218),
    .X(_3395_));
 sky130_fd_sc_hd__o2111a_1 _6249_ (.A1(net211),
    .A2(_3082_),
    .B1(_3392_),
    .C1(_3393_),
    .D1(_3395_),
    .X(_3396_));
 sky130_fd_sc_hd__o21ai_1 _6250_ (.A1(net282),
    .A2(_3386_),
    .B1(_3396_),
    .Y(_3397_));
 sky130_fd_sc_hd__a21o_1 _6251_ (.A1(_1601_),
    .A2(_1603_),
    .B1(net218),
    .X(_3398_));
 sky130_fd_sc_hd__and3_1 _6252_ (.A(net429),
    .B(_3397_),
    .C(_3398_),
    .X(_0654_));
 sky130_fd_sc_hd__a21boi_2 _6253_ (.A1(_3382_),
    .A2(_3385_),
    .B1_N(_3383_),
    .Y(_3399_));
 sky130_fd_sc_hd__xnor2_1 _6254_ (.A(_1591_),
    .B(net313),
    .Y(_3400_));
 sky130_fd_sc_hd__nor2_1 _6255_ (.A(_1594_),
    .B(_3400_),
    .Y(_3401_));
 sky130_fd_sc_hd__nand2_1 _6256_ (.A(_1594_),
    .B(_3400_),
    .Y(_3402_));
 sky130_fd_sc_hd__nand2b_1 _6257_ (.A_N(_3401_),
    .B(_3402_),
    .Y(_3403_));
 sky130_fd_sc_hd__xnor2_1 _6258_ (.A(_3399_),
    .B(_3403_),
    .Y(_3404_));
 sky130_fd_sc_hd__mux4_1 _6259_ (.A0(_1594_),
    .A1(_1603_),
    .A2(_1656_),
    .A3(_1627_),
    .S0(net191),
    .S1(net202),
    .X(_3405_));
 sky130_fd_sc_hd__mux2_1 _6260_ (.A0(_3337_),
    .A1(_3405_),
    .S(net199),
    .X(_3406_));
 sky130_fd_sc_hd__mux2_1 _6261_ (.A0(_3267_),
    .A1(_3406_),
    .S(net207),
    .X(_3407_));
 sky130_fd_sc_hd__nand2_1 _6262_ (.A(net211),
    .B(_3106_),
    .Y(_3408_));
 sky130_fd_sc_hd__o211a_1 _6263_ (.A1(net211),
    .A2(_3407_),
    .B1(_3408_),
    .C1(_2720_),
    .X(_3409_));
 sky130_fd_sc_hd__o21ai_1 _6264_ (.A1(net211),
    .A2(_3112_),
    .B1(_3126_),
    .Y(_3410_));
 sky130_fd_sc_hd__a21o_1 _6265_ (.A1(_1594_),
    .A2(net310),
    .B1(_1591_),
    .X(_3411_));
 sky130_fd_sc_hd__a221oi_1 _6266_ (.A1(_1595_),
    .A2(_2713_),
    .B1(net281),
    .B2(_3411_),
    .C1(net220),
    .Y(_3412_));
 sky130_fd_sc_hd__o311a_1 _6267_ (.A1(net211),
    .A2(_2922_),
    .A3(_2923_),
    .B1(_3410_),
    .C1(_3412_),
    .X(_3413_));
 sky130_fd_sc_hd__o21ai_1 _6268_ (.A1(net282),
    .A2(_3404_),
    .B1(_3413_),
    .Y(_3414_));
 sky130_fd_sc_hd__a21o_1 _6269_ (.A1(_1591_),
    .A2(_1594_),
    .B1(net218),
    .X(_3415_));
 sky130_fd_sc_hd__o211a_1 _6270_ (.A1(_3409_),
    .A2(_3414_),
    .B1(_3415_),
    .C1(net435),
    .X(_0655_));
 sky130_fd_sc_hd__o21ai_1 _6271_ (.A1(_3399_),
    .A2(_3401_),
    .B1(_3402_),
    .Y(_3416_));
 sky130_fd_sc_hd__or2_1 _6272_ (.A(_1641_),
    .B(net316),
    .X(_3417_));
 sky130_fd_sc_hd__nand2_1 _6273_ (.A(_1641_),
    .B(net316),
    .Y(_3418_));
 sky130_fd_sc_hd__nand2_1 _6274_ (.A(_1641_),
    .B(net313),
    .Y(_3419_));
 sky130_fd_sc_hd__or2_1 _6275_ (.A(_1641_),
    .B(net313),
    .X(_3420_));
 sky130_fd_sc_hd__o2111a_1 _6276_ (.A1(_3399_),
    .A2(_3401_),
    .B1(_3402_),
    .C1(_3419_),
    .D1(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__a311o_1 _6277_ (.A1(_3416_),
    .A2(_3417_),
    .A3(_3418_),
    .B1(_3421_),
    .C1(net282),
    .X(_3422_));
 sky130_fd_sc_hd__a31o_1 _6278_ (.A1(net205),
    .A2(net192),
    .A3(_1594_),
    .B1(_2830_),
    .X(_3423_));
 sky130_fd_sc_hd__a211o_1 _6279_ (.A1(net202),
    .A2(_3387_),
    .B1(_3423_),
    .C1(net196),
    .X(_3424_));
 sky130_fd_sc_hd__o211a_1 _6280_ (.A1(net199),
    .A2(_3355_),
    .B1(_3424_),
    .C1(net208),
    .X(_3425_));
 sky130_fd_sc_hd__a211o_1 _6281_ (.A1(net186),
    .A2(_3286_),
    .B1(_3425_),
    .C1(net212),
    .X(_3426_));
 sky130_fd_sc_hd__o211a_1 _6282_ (.A1(net216),
    .A2(_3133_),
    .B1(_3426_),
    .C1(_2720_),
    .X(_3427_));
 sky130_fd_sc_hd__a221o_1 _6283_ (.A1(_1638_),
    .A2(_2671_),
    .B1(_2717_),
    .B2(_1635_),
    .C1(net220),
    .X(_3428_));
 sky130_fd_sc_hd__a221o_1 _6284_ (.A1(_1641_),
    .A2(_2713_),
    .B1(net310),
    .B2(_1639_),
    .C1(_3428_),
    .X(_3429_));
 sky130_fd_sc_hd__a211oi_1 _6285_ (.A1(_3128_),
    .A2(_3136_),
    .B1(_3427_),
    .C1(_3429_),
    .Y(_3430_));
 sky130_fd_sc_hd__a221oi_2 _6286_ (.A1(net2298),
    .A2(net220),
    .B1(_3422_),
    .B2(_3430_),
    .C1(net63),
    .Y(_0656_));
 sky130_fd_sc_hd__and2_1 _6287_ (.A(net453),
    .B(net642),
    .X(_0657_));
 sky130_fd_sc_hd__and2_1 _6288_ (.A(net451),
    .B(net666),
    .X(_0658_));
 sky130_fd_sc_hd__and2_1 _6289_ (.A(net450),
    .B(net596),
    .X(_0659_));
 sky130_fd_sc_hd__and2_1 _6290_ (.A(net449),
    .B(net604),
    .X(_0660_));
 sky130_fd_sc_hd__and2_1 _6291_ (.A(net448),
    .B(net575),
    .X(_0661_));
 sky130_fd_sc_hd__and2_1 _6292_ (.A(net442),
    .B(net634),
    .X(_0662_));
 sky130_fd_sc_hd__and2_1 _6293_ (.A(net442),
    .B(net613),
    .X(_0663_));
 sky130_fd_sc_hd__and2_1 _6294_ (.A(net450),
    .B(net585),
    .X(_0664_));
 sky130_fd_sc_hd__and2_1 _6295_ (.A(net435),
    .B(net617),
    .X(_0665_));
 sky130_fd_sc_hd__and2_1 _6296_ (.A(net429),
    .B(net732),
    .X(_0666_));
 sky130_fd_sc_hd__and2_1 _6297_ (.A(net449),
    .B(net674),
    .X(_0667_));
 sky130_fd_sc_hd__and2_1 _6298_ (.A(net443),
    .B(net567),
    .X(_0668_));
 sky130_fd_sc_hd__and2_1 _6299_ (.A(net449),
    .B(net646),
    .X(_0669_));
 sky130_fd_sc_hd__and2_1 _6300_ (.A(net442),
    .B(net692),
    .X(_0670_));
 sky130_fd_sc_hd__and2_1 _6301_ (.A(net443),
    .B(net650),
    .X(_0671_));
 sky130_fd_sc_hd__and2_1 _6302_ (.A(net443),
    .B(net543),
    .X(_0672_));
 sky130_fd_sc_hd__and2_1 _6303_ (.A(net454),
    .B(net771),
    .X(_0673_));
 sky130_fd_sc_hd__and2_1 _6304_ (.A(net438),
    .B(net694),
    .X(_0674_));
 sky130_fd_sc_hd__and2_1 _6305_ (.A(net432),
    .B(net684),
    .X(_0675_));
 sky130_fd_sc_hd__and2_1 _6306_ (.A(net431),
    .B(net581),
    .X(_0676_));
 sky130_fd_sc_hd__and2_1 _6307_ (.A(net430),
    .B(net630),
    .X(_0677_));
 sky130_fd_sc_hd__and2_1 _6308_ (.A(net432),
    .B(net682),
    .X(_0678_));
 sky130_fd_sc_hd__and2_1 _6309_ (.A(net436),
    .B(net782),
    .X(_0679_));
 sky130_fd_sc_hd__and2_1 _6310_ (.A(net432),
    .B(net752),
    .X(_0680_));
 sky130_fd_sc_hd__and2_1 _6311_ (.A(net431),
    .B(net658),
    .X(_0681_));
 sky130_fd_sc_hd__and2_1 _6312_ (.A(net431),
    .B(net696),
    .X(_0682_));
 sky130_fd_sc_hd__and2_1 _6313_ (.A(net430),
    .B(net557),
    .X(_0683_));
 sky130_fd_sc_hd__and2_1 _6314_ (.A(net429),
    .B(net776),
    .X(_0684_));
 sky130_fd_sc_hd__and2_1 _6315_ (.A(net429),
    .B(net594),
    .X(_0685_));
 sky130_fd_sc_hd__and2_1 _6316_ (.A(net431),
    .B(net726),
    .X(_0686_));
 sky130_fd_sc_hd__and2_1 _6317_ (.A(net2006),
    .B(net453),
    .X(_0687_));
 sky130_fd_sc_hd__and2_1 _6318_ (.A(net2059),
    .B(net453),
    .X(_0688_));
 sky130_fd_sc_hd__and2_1 _6319_ (.A(net1308),
    .B(net453),
    .X(_0689_));
 sky130_fd_sc_hd__and2_1 _6320_ (.A(net1631),
    .B(net453),
    .X(_0690_));
 sky130_fd_sc_hd__and2_1 _6321_ (.A(_2620_),
    .B(net320),
    .X(_3431_));
 sky130_fd_sc_hd__nand2_1 _6322_ (.A(_2620_),
    .B(net320),
    .Y(_3432_));
 sky130_fd_sc_hd__nor2_1 _6323_ (.A(net460),
    .B(net280),
    .Y(_3433_));
 sky130_fd_sc_hd__nand2_1 _6324_ (.A(net447),
    .B(_3432_),
    .Y(_3434_));
 sky130_fd_sc_hd__o22a_1 _6325_ (.A1(net298),
    .A2(_3432_),
    .B1(_3434_),
    .B2(net885),
    .X(_0691_));
 sky130_fd_sc_hd__o22a_1 _6326_ (.A1(net299),
    .A2(_3432_),
    .B1(_3434_),
    .B2(net1063),
    .X(_0692_));
 sky130_fd_sc_hd__o22a_1 _6327_ (.A1(net353),
    .A2(_3432_),
    .B1(_3434_),
    .B2(net907),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _6328_ (.A1(net355),
    .A2(net280),
    .B1(net233),
    .B2(net979),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _6329_ (.A1(net356),
    .A2(net280),
    .B1(net233),
    .B2(net1697),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _6330_ (.A1(net354),
    .A2(net280),
    .B1(net233),
    .B2(net1266),
    .X(_0696_));
 sky130_fd_sc_hd__a22o_1 _6331_ (.A1(net352),
    .A2(net279),
    .B1(net232),
    .B2(net1477),
    .X(_0697_));
 sky130_fd_sc_hd__a22o_1 _6332_ (.A1(net351),
    .A2(net280),
    .B1(net233),
    .B2(net1329),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _6333_ (.A1(net358),
    .A2(net279),
    .B1(net232),
    .B2(net1591),
    .X(_0699_));
 sky130_fd_sc_hd__a22o_1 _6334_ (.A1(net359),
    .A2(net280),
    .B1(net233),
    .B2(net1272),
    .X(_0700_));
 sky130_fd_sc_hd__a22o_1 _6335_ (.A1(net357),
    .A2(net279),
    .B1(net232),
    .B2(net1302),
    .X(_0701_));
 sky130_fd_sc_hd__a22o_1 _6336_ (.A1(net361),
    .A2(net279),
    .B1(net232),
    .B2(net1672),
    .X(_0702_));
 sky130_fd_sc_hd__a22o_1 _6337_ (.A1(_1349_),
    .A2(net280),
    .B1(net233),
    .B2(net1089),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _6338_ (.A1(net360),
    .A2(net279),
    .B1(net232),
    .B2(net1413),
    .X(_0704_));
 sky130_fd_sc_hd__a22o_1 _6339_ (.A1(net350),
    .A2(net280),
    .B1(net233),
    .B2(net1278),
    .X(_0705_));
 sky130_fd_sc_hd__a22o_1 _6340_ (.A1(net349),
    .A2(net280),
    .B1(net233),
    .B2(net1515),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _6341_ (.A1(net345),
    .A2(net280),
    .B1(net233),
    .B2(net1451),
    .X(_0707_));
 sky130_fd_sc_hd__a22o_1 _6342_ (.A1(net344),
    .A2(net280),
    .B1(net233),
    .B2(net1627),
    .X(_0708_));
 sky130_fd_sc_hd__a22o_1 _6343_ (.A1(net341),
    .A2(net280),
    .B1(net233),
    .B2(net1756),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _6344_ (.A1(net343),
    .A2(net279),
    .B1(net232),
    .B2(net1316),
    .X(_0710_));
 sky130_fd_sc_hd__a22o_1 _6345_ (.A1(net342),
    .A2(net279),
    .B1(net232),
    .B2(net1208),
    .X(_0711_));
 sky130_fd_sc_hd__a22o_1 _6346_ (.A1(net346),
    .A2(net279),
    .B1(net232),
    .B2(net1521),
    .X(_0712_));
 sky130_fd_sc_hd__a22o_1 _6347_ (.A1(net348),
    .A2(net280),
    .B1(net233),
    .B2(net1779),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _6348_ (.A1(net347),
    .A2(net279),
    .B1(net232),
    .B2(net999),
    .X(_0714_));
 sky130_fd_sc_hd__a22o_1 _6349_ (.A1(net334),
    .A2(net280),
    .B1(net233),
    .B2(net1224),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _6350_ (.A1(net337),
    .A2(net279),
    .B1(net232),
    .B2(net1373),
    .X(_0716_));
 sky130_fd_sc_hd__a22o_1 _6351_ (.A1(net338),
    .A2(net279),
    .B1(net232),
    .B2(net1491),
    .X(_0717_));
 sky130_fd_sc_hd__a22o_1 _6352_ (.A1(net336),
    .A2(net279),
    .B1(net232),
    .B2(net1055),
    .X(_0718_));
 sky130_fd_sc_hd__a22o_1 _6353_ (.A1(net333),
    .A2(net279),
    .B1(net232),
    .B2(net993),
    .X(_0719_));
 sky130_fd_sc_hd__a22o_1 _6354_ (.A1(net339),
    .A2(net279),
    .B1(net232),
    .B2(net1537),
    .X(_0720_));
 sky130_fd_sc_hd__a22o_1 _6355_ (.A1(net340),
    .A2(net279),
    .B1(net232),
    .B2(net1375),
    .X(_0721_));
 sky130_fd_sc_hd__a22o_1 _6356_ (.A1(net335),
    .A2(net279),
    .B1(net232),
    .B2(net1569),
    .X(_0722_));
 sky130_fd_sc_hd__nor2_2 _6357_ (.A(_2509_),
    .B(_2580_),
    .Y(_3435_));
 sky130_fd_sc_hd__or2_1 _6358_ (.A(_2509_),
    .B(_2580_),
    .X(_3436_));
 sky130_fd_sc_hd__nor2_1 _6359_ (.A(net460),
    .B(net278),
    .Y(_3437_));
 sky130_fd_sc_hd__nand2_1 _6360_ (.A(net454),
    .B(_3436_),
    .Y(_3438_));
 sky130_fd_sc_hd__o22a_1 _6361_ (.A1(net298),
    .A2(_3436_),
    .B1(_3438_),
    .B2(net931),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _6362_ (.A1(net299),
    .A2(net278),
    .B1(net231),
    .B2(net1343),
    .X(_0724_));
 sky130_fd_sc_hd__a22o_1 _6363_ (.A1(_1462_),
    .A2(net278),
    .B1(net231),
    .B2(net1220),
    .X(_0725_));
 sky130_fd_sc_hd__o22a_1 _6364_ (.A1(net355),
    .A2(_3436_),
    .B1(_3438_),
    .B2(net909),
    .X(_0726_));
 sky130_fd_sc_hd__a22o_1 _6365_ (.A1(net356),
    .A2(net278),
    .B1(net231),
    .B2(net1750),
    .X(_0727_));
 sky130_fd_sc_hd__a22o_1 _6366_ (.A1(net354),
    .A2(net278),
    .B1(net231),
    .B2(net1517),
    .X(_0728_));
 sky130_fd_sc_hd__a22o_1 _6367_ (.A1(net352),
    .A2(net277),
    .B1(net230),
    .B2(net1365),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _6368_ (.A1(net351),
    .A2(net278),
    .B1(net231),
    .B2(net1647),
    .X(_0730_));
 sky130_fd_sc_hd__a22o_1 _6369_ (.A1(net358),
    .A2(net278),
    .B1(net231),
    .B2(net1357),
    .X(_0731_));
 sky130_fd_sc_hd__a22o_1 _6370_ (.A1(net359),
    .A2(net278),
    .B1(net231),
    .B2(net967),
    .X(_0732_));
 sky130_fd_sc_hd__a22o_1 _6371_ (.A1(net357),
    .A2(net277),
    .B1(net230),
    .B2(net1135),
    .X(_0733_));
 sky130_fd_sc_hd__a22o_1 _6372_ (.A1(net361),
    .A2(net277),
    .B1(net230),
    .B2(net1337),
    .X(_0734_));
 sky130_fd_sc_hd__a22o_1 _6373_ (.A1(_1349_),
    .A2(net278),
    .B1(net231),
    .B2(net1280),
    .X(_0735_));
 sky130_fd_sc_hd__a22o_1 _6374_ (.A1(net360),
    .A2(net277),
    .B1(net230),
    .B2(net1409),
    .X(_0736_));
 sky130_fd_sc_hd__a22o_1 _6375_ (.A1(net350),
    .A2(net278),
    .B1(net231),
    .B2(net1603),
    .X(_0737_));
 sky130_fd_sc_hd__a22o_1 _6376_ (.A1(net349),
    .A2(net278),
    .B1(net231),
    .B2(net1085),
    .X(_0738_));
 sky130_fd_sc_hd__a22o_1 _6377_ (.A1(net345),
    .A2(net277),
    .B1(net230),
    .B2(net1127),
    .X(_0739_));
 sky130_fd_sc_hd__a22o_1 _6378_ (.A1(net344),
    .A2(net278),
    .B1(net231),
    .B2(net1417),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _6379_ (.A1(net341),
    .A2(net278),
    .B1(net231),
    .B2(net1359),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _6380_ (.A1(net343),
    .A2(net277),
    .B1(net230),
    .B2(net1519),
    .X(_0742_));
 sky130_fd_sc_hd__a22o_1 _6381_ (.A1(net342),
    .A2(net277),
    .B1(net230),
    .B2(net1250),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _6382_ (.A1(net346),
    .A2(net277),
    .B1(net230),
    .B2(net1115),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _6383_ (.A1(net348),
    .A2(net278),
    .B1(net231),
    .B2(net1314),
    .X(_0745_));
 sky130_fd_sc_hd__a22o_1 _6384_ (.A1(net347),
    .A2(net277),
    .B1(net230),
    .B2(net1443),
    .X(_0746_));
 sky130_fd_sc_hd__a22o_1 _6385_ (.A1(net334),
    .A2(net278),
    .B1(net231),
    .B2(net1333),
    .X(_0747_));
 sky130_fd_sc_hd__a22o_1 _6386_ (.A1(net337),
    .A2(net277),
    .B1(net230),
    .B2(net1509),
    .X(_0748_));
 sky130_fd_sc_hd__a22o_1 _6387_ (.A1(net338),
    .A2(net277),
    .B1(net230),
    .B2(net1465),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _6388_ (.A1(net336),
    .A2(net277),
    .B1(net230),
    .B2(net1369),
    .X(_0750_));
 sky130_fd_sc_hd__a22o_1 _6389_ (.A1(_1651_),
    .A2(net277),
    .B1(net230),
    .B2(net1200),
    .X(_0751_));
 sky130_fd_sc_hd__a22o_1 _6390_ (.A1(net339),
    .A2(net277),
    .B1(net230),
    .B2(net1914),
    .X(_0752_));
 sky130_fd_sc_hd__a22o_1 _6391_ (.A1(net340),
    .A2(net277),
    .B1(net230),
    .B2(net1226),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _6392_ (.A1(net335),
    .A2(net277),
    .B1(net230),
    .B2(net1686),
    .X(_0754_));
 sky130_fd_sc_hd__a21o_1 _6393_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .A2(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .B1(net773),
    .X(_3439_));
 sky130_fd_sc_hd__and3_1 _6394_ (.A(net448),
    .B(_1822_),
    .C(net774),
    .X(_0755_));
 sky130_fd_sc_hd__or2_1 _6395_ (.A(net464),
    .B(_1823_),
    .X(_3440_));
 sky130_fd_sc_hd__a21oi_1 _6396_ (.A1(net828),
    .A2(_1822_),
    .B1(_3440_),
    .Y(_0756_));
 sky130_fd_sc_hd__nor2_1 _6397_ (.A(net464),
    .B(net2285),
    .Y(_0757_));
 sky130_fd_sc_hd__nor2_1 _6398_ (.A(net463),
    .B(net2110),
    .Y(_0758_));
 sky130_fd_sc_hd__and2_1 _6399_ (.A(net450),
    .B(net2277),
    .X(_0759_));
 sky130_fd_sc_hd__and2_1 _6400_ (.A(net449),
    .B(net2070),
    .X(_0760_));
 sky130_fd_sc_hd__and2_1 _6401_ (.A(net448),
    .B(net2236),
    .X(_0761_));
 sky130_fd_sc_hd__and2_1 _6402_ (.A(net442),
    .B(net2191),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _6403_ (.A(net460),
    .B(net2141),
    .Y(_0763_));
 sky130_fd_sc_hd__and2_1 _6404_ (.A(net450),
    .B(_1935_),
    .X(_0764_));
 sky130_fd_sc_hd__and2_1 _6405_ (.A(net440),
    .B(net2216),
    .X(_0765_));
 sky130_fd_sc_hd__nor2_1 _6406_ (.A(net457),
    .B(net2214),
    .Y(_0766_));
 sky130_fd_sc_hd__and2_1 _6407_ (.A(net449),
    .B(net2099),
    .X(_0767_));
 sky130_fd_sc_hd__and2_1 _6408_ (.A(net442),
    .B(net2172),
    .X(_0768_));
 sky130_fd_sc_hd__nor2_1 _6409_ (.A(net461),
    .B(net2271),
    .Y(_0769_));
 sky130_fd_sc_hd__and2_1 _6410_ (.A(net442),
    .B(net2091),
    .X(_0770_));
 sky130_fd_sc_hd__and2_1 _6411_ (.A(net443),
    .B(net2244),
    .X(_0771_));
 sky130_fd_sc_hd__and2_1 _6412_ (.A(net443),
    .B(net2137),
    .X(_0772_));
 sky130_fd_sc_hd__and2_1 _6413_ (.A(net453),
    .B(net2200),
    .X(_0773_));
 sky130_fd_sc_hd__and2_1 _6414_ (.A(net438),
    .B(_1913_),
    .X(_0774_));
 sky130_fd_sc_hd__nor2_1 _6415_ (.A(net459),
    .B(net2123),
    .Y(_0775_));
 sky130_fd_sc_hd__and2_1 _6416_ (.A(net432),
    .B(net2080),
    .X(_0776_));
 sky130_fd_sc_hd__and2_1 _6417_ (.A(net430),
    .B(net2154),
    .X(_0777_));
 sky130_fd_sc_hd__nor2_1 _6418_ (.A(net458),
    .B(net2180),
    .Y(_0778_));
 sky130_fd_sc_hd__and2_1 _6419_ (.A(net432),
    .B(net2241),
    .X(_0779_));
 sky130_fd_sc_hd__nor2_1 _6420_ (.A(net458),
    .B(net2116),
    .Y(_0780_));
 sky130_fd_sc_hd__nor2_1 _6421_ (.A(net458),
    .B(net2158),
    .Y(_0781_));
 sky130_fd_sc_hd__nor2_1 _6422_ (.A(net458),
    .B(_1891_),
    .Y(_0782_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(net457),
    .B(_1888_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor2_1 _6424_ (.A(net457),
    .B(net2185),
    .Y(_0784_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(net429),
    .B(net2176),
    .X(_0785_));
 sky130_fd_sc_hd__and2_1 _6426_ (.A(net431),
    .B(net2229),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_1 _6427_ (.A(_2035_),
    .B(net162),
    .Y(_0787_));
 sky130_fd_sc_hd__nor2_1 _6428_ (.A(net162),
    .B(_2477_),
    .Y(_0788_));
 sky130_fd_sc_hd__and3_1 _6429_ (.A(_1282_),
    .B(_2034_),
    .C(net175),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(net1959),
    .B(net179),
    .X(_0790_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(net1946),
    .B(net182),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(net2042),
    .B(net180),
    .X(_0792_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(net608),
    .B(net180),
    .X(_0793_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ),
    .B(net180),
    .X(_0794_));
 sky130_fd_sc_hd__and2_1 _6435_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ),
    .B(net177),
    .X(_0795_));
 sky130_fd_sc_hd__and2_1 _6436_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ),
    .B(net180),
    .X(_0796_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ),
    .B(net179),
    .X(_0797_));
 sky130_fd_sc_hd__and2_1 _6438_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ),
    .B(net178),
    .X(_0798_));
 sky130_fd_sc_hd__and2_1 _6439_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ),
    .B(net178),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ),
    .B(net177),
    .X(_0800_));
 sky130_fd_sc_hd__and2_1 _6441_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ),
    .B(net177),
    .X(_0801_));
 sky130_fd_sc_hd__and2_1 _6442_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ),
    .B(net177),
    .X(_0802_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ),
    .B(net179),
    .X(_0803_));
 sky130_fd_sc_hd__and2_1 _6444_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ),
    .B(net177),
    .X(_0804_));
 sky130_fd_sc_hd__and2_1 _6445_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ),
    .B(net172),
    .X(_0805_));
 sky130_fd_sc_hd__and2_1 _6446_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ),
    .B(net178),
    .X(_0806_));
 sky130_fd_sc_hd__and2_1 _6447_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ),
    .B(net173),
    .X(_0807_));
 sky130_fd_sc_hd__and2_1 _6448_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ),
    .B(net178),
    .X(_0808_));
 sky130_fd_sc_hd__and2_1 _6449_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ),
    .B(net179),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _6450_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ),
    .B(net177),
    .X(_0810_));
 sky130_fd_sc_hd__and2_1 _6451_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ),
    .B(net180),
    .X(_0811_));
 sky130_fd_sc_hd__and2_1 _6452_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ),
    .B(net180),
    .X(_0812_));
 sky130_fd_sc_hd__and2_1 _6453_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ),
    .B(net173),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _6454_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ),
    .B(net173),
    .X(_0814_));
 sky130_fd_sc_hd__and2_1 _6455_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ),
    .B(net173),
    .X(_0815_));
 sky130_fd_sc_hd__and2_1 _6456_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ),
    .B(net173),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _6457_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ),
    .B(net174),
    .X(_0817_));
 sky130_fd_sc_hd__and2_1 _6458_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ),
    .B(net180),
    .X(_0818_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ),
    .B(net174),
    .X(_0819_));
 sky130_fd_sc_hd__and2_1 _6460_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ),
    .B(net174),
    .X(_0820_));
 sky130_fd_sc_hd__and2_1 _6461_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ),
    .B(net174),
    .X(_0821_));
 sky130_fd_sc_hd__and2_1 _6462_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ),
    .B(net172),
    .X(_0822_));
 sky130_fd_sc_hd__and2_1 _6463_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ),
    .B(net172),
    .X(_0823_));
 sky130_fd_sc_hd__and2_1 _6464_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ),
    .B(net173),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _6465_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ),
    .B(net173),
    .X(_0825_));
 sky130_fd_sc_hd__and2_1 _6466_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ),
    .B(net177),
    .X(_0826_));
 sky130_fd_sc_hd__and2_1 _6467_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ),
    .B(net177),
    .X(_0827_));
 sky130_fd_sc_hd__and2_1 _6468_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ),
    .B(net180),
    .X(_0828_));
 sky130_fd_sc_hd__and2_1 _6469_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ),
    .B(net181),
    .X(_0829_));
 sky130_fd_sc_hd__and2_1 _6470_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ),
    .B(net180),
    .X(_0830_));
 sky130_fd_sc_hd__and2_1 _6471_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ),
    .B(net178),
    .X(_0831_));
 sky130_fd_sc_hd__and2_1 _6472_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ),
    .B(net177),
    .X(_0832_));
 sky130_fd_sc_hd__and2_1 _6473_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ),
    .B(net182),
    .X(_0833_));
 sky130_fd_sc_hd__and2_1 _6474_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ),
    .B(net177),
    .X(_0834_));
 sky130_fd_sc_hd__and2_1 _6475_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ),
    .B(net178),
    .X(_0835_));
 sky130_fd_sc_hd__and2_1 _6476_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ),
    .B(net177),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _6477_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ),
    .B(net172),
    .X(_0837_));
 sky130_fd_sc_hd__and2_1 _6478_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ),
    .B(net178),
    .X(_0838_));
 sky130_fd_sc_hd__and2_1 _6479_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ),
    .B(net174),
    .X(_0839_));
 sky130_fd_sc_hd__and2_1 _6480_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ),
    .B(net179),
    .X(_0840_));
 sky130_fd_sc_hd__and2_1 _6481_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ),
    .B(net179),
    .X(_0841_));
 sky130_fd_sc_hd__and2_1 _6482_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ),
    .B(net177),
    .X(_0842_));
 sky130_fd_sc_hd__and2_1 _6483_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ),
    .B(net177),
    .X(_0843_));
 sky130_fd_sc_hd__and2_1 _6484_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ),
    .B(net180),
    .X(_0844_));
 sky130_fd_sc_hd__and2_1 _6485_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ),
    .B(net173),
    .X(_0845_));
 sky130_fd_sc_hd__and2_1 _6486_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ),
    .B(net173),
    .X(_0846_));
 sky130_fd_sc_hd__and2_1 _6487_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ),
    .B(net173),
    .X(_0847_));
 sky130_fd_sc_hd__and2_1 _6488_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ),
    .B(net177),
    .X(_0848_));
 sky130_fd_sc_hd__and2_1 _6489_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ),
    .B(net174),
    .X(_0849_));
 sky130_fd_sc_hd__and2_1 _6490_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ),
    .B(net180),
    .X(_0850_));
 sky130_fd_sc_hd__and2_1 _6491_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ),
    .B(net173),
    .X(_0851_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ),
    .B(net174),
    .X(_0852_));
 sky130_fd_sc_hd__and2_1 _6493_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ),
    .B(net173),
    .X(_0853_));
 sky130_fd_sc_hd__and2_1 _6494_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ),
    .B(net172),
    .X(_0854_));
 sky130_fd_sc_hd__and2_1 _6495_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ),
    .B(net172),
    .X(_0855_));
 sky130_fd_sc_hd__and2_1 _6496_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ),
    .B(net173),
    .X(_0856_));
 sky130_fd_sc_hd__and2_1 _6497_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ),
    .B(net173),
    .X(_0857_));
 sky130_fd_sc_hd__and2_1 _6498_ (.A(net424),
    .B(net181),
    .X(_0858_));
 sky130_fd_sc_hd__and2_1 _6499_ (.A(net414),
    .B(net181),
    .X(_0859_));
 sky130_fd_sc_hd__and2_1 _6500_ (.A(net403),
    .B(net180),
    .X(_0860_));
 sky130_fd_sc_hd__and2_1 _6501_ (.A(net2126),
    .B(net180),
    .X(_0861_));
 sky130_fd_sc_hd__and2_1 _6502_ (.A(net395),
    .B(net181),
    .X(_0862_));
 sky130_fd_sc_hd__and2_1 _6503_ (.A(net385),
    .B(net181),
    .X(_0863_));
 sky130_fd_sc_hd__and2_1 _6504_ (.A(net374),
    .B(net181),
    .X(_0864_));
 sky130_fd_sc_hd__and2_1 _6505_ (.A(net369),
    .B(net180),
    .X(_0865_));
 sky130_fd_sc_hd__and2_1 _6506_ (.A(net822),
    .B(net182),
    .X(_0866_));
 sky130_fd_sc_hd__and2_1 _6507_ (.A(net769),
    .B(net179),
    .X(_0867_));
 sky130_fd_sc_hd__and2_1 _6508_ (.A(net849),
    .B(net179),
    .X(_0868_));
 sky130_fd_sc_hd__and2_1 _6509_ (.A(net812),
    .B(net178),
    .X(_0869_));
 sky130_fd_sc_hd__and2_1 _6510_ (.A(net841),
    .B(net177),
    .X(_0870_));
 sky130_fd_sc_hd__and2_1 _6511_ (.A(net796),
    .B(net175),
    .X(_0871_));
 sky130_fd_sc_hd__and2_1 _6512_ (.A(net865),
    .B(net175),
    .X(_0872_));
 sky130_fd_sc_hd__and2_1 _6513_ (.A(net804),
    .B(net178),
    .X(_0873_));
 sky130_fd_sc_hd__and2_1 _6514_ (.A(net1010),
    .B(net174),
    .X(_0874_));
 sky130_fd_sc_hd__and2_1 _6515_ (.A(net887),
    .B(net179),
    .X(_0875_));
 sky130_fd_sc_hd__and2_1 _6516_ (.A(net843),
    .B(net178),
    .X(_0876_));
 sky130_fd_sc_hd__and2_1 _6517_ (.A(net561),
    .B(net177),
    .X(_0877_));
 sky130_fd_sc_hd__and2_1 _6518_ (.A(net832),
    .B(net178),
    .X(_0878_));
 sky130_fd_sc_hd__and2_1 _6519_ (.A(net571),
    .B(net179),
    .X(_0879_));
 sky130_fd_sc_hd__and2_1 _6520_ (.A(net541),
    .B(net182),
    .X(_0880_));
 sky130_fd_sc_hd__and2_1 _6521_ (.A(net791),
    .B(net182),
    .X(_0881_));
 sky130_fd_sc_hd__and2_1 _6522_ (.A(net609),
    .B(net178),
    .X(_0882_));
 sky130_fd_sc_hd__and2_1 _6523_ (.A(net835),
    .B(net173),
    .X(_0883_));
 sky130_fd_sc_hd__and2_1 _6524_ (.A(net891),
    .B(net171),
    .X(_0884_));
 sky130_fd_sc_hd__and2_1 _6525_ (.A(net869),
    .B(net171),
    .X(_0885_));
 sky130_fd_sc_hd__and2_1 _6526_ (.A(net845),
    .B(net171),
    .X(_0886_));
 sky130_fd_sc_hd__and2_1 _6527_ (.A(net897),
    .B(net171),
    .X(_0887_));
 sky130_fd_sc_hd__and2_1 _6528_ (.A(net974),
    .B(net171),
    .X(_0888_));
 sky130_fd_sc_hd__and2_1 _6529_ (.A(net816),
    .B(net171),
    .X(_0889_));
 sky130_fd_sc_hd__and2_1 _6530_ (.A(net883),
    .B(net171),
    .X(_0890_));
 sky130_fd_sc_hd__and2_1 _6531_ (.A(net644),
    .B(net171),
    .X(_0891_));
 sky130_fd_sc_hd__and2_1 _6532_ (.A(net879),
    .B(net172),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _6533_ (.A(net563),
    .B(net172),
    .X(_0893_));
 sky130_fd_sc_hd__and2_1 _6534_ (.A(net800),
    .B(net172),
    .X(_0894_));
 sky130_fd_sc_hd__and2_1 _6535_ (.A(net818),
    .B(net172),
    .X(_0895_));
 sky130_fd_sc_hd__and2_1 _6536_ (.A(net873),
    .B(net180),
    .X(_0896_));
 sky130_fd_sc_hd__and2_1 _6537_ (.A(net839),
    .B(net178),
    .X(_0897_));
 sky130_fd_sc_hd__and2_1 _6538_ (.A(net628),
    .B(net178),
    .X(_0898_));
 sky130_fd_sc_hd__and2_1 _6539_ (.A(net606),
    .B(net179),
    .X(_0899_));
 sky130_fd_sc_hd__and2_1 _6540_ (.A(net551),
    .B(net176),
    .X(_0900_));
 sky130_fd_sc_hd__and2_1 _6541_ (.A(net875),
    .B(net175),
    .X(_0901_));
 sky130_fd_sc_hd__and2_1 _6542_ (.A(net778),
    .B(net175),
    .X(_0902_));
 sky130_fd_sc_hd__and2_1 _6543_ (.A(net814),
    .B(net178),
    .X(_0903_));
 sky130_fd_sc_hd__and2_1 _6544_ (.A(net754),
    .B(net174),
    .X(_0904_));
 sky130_fd_sc_hd__and2_1 _6545_ (.A(net539),
    .B(net172),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _6546_ (.A(net830),
    .B(net178),
    .X(_0906_));
 sky130_fd_sc_hd__and2_1 _6547_ (.A(net559),
    .B(net176),
    .X(_0907_));
 sky130_fd_sc_hd__and2_1 _6548_ (.A(net847),
    .B(net179),
    .X(_0908_));
 sky130_fd_sc_hd__and2_1 _6549_ (.A(net856),
    .B(net179),
    .X(_0909_));
 sky130_fd_sc_hd__and2_1 _6550_ (.A(net802),
    .B(net176),
    .X(_0910_));
 sky130_fd_sc_hd__and2_1 _6551_ (.A(net793),
    .B(net180),
    .X(_0911_));
 sky130_fd_sc_hd__and2_1 _6552_ (.A(net758),
    .B(net181),
    .X(_0912_));
 sky130_fd_sc_hd__and2_1 _6553_ (.A(net718),
    .B(net173),
    .X(_0913_));
 sky130_fd_sc_hd__and2_1 _6554_ (.A(net810),
    .B(net171),
    .X(_0914_));
 sky130_fd_sc_hd__and2_1 _6555_ (.A(net656),
    .B(net171),
    .X(_0915_));
 sky130_fd_sc_hd__and2_1 _6556_ (.A(net863),
    .B(net172),
    .X(_0916_));
 sky130_fd_sc_hd__and2_1 _6557_ (.A(net861),
    .B(net171),
    .X(_0917_));
 sky130_fd_sc_hd__and2_1 _6558_ (.A(net2053),
    .B(net171),
    .X(_0918_));
 sky130_fd_sc_hd__and2_1 _6559_ (.A(net824),
    .B(net171),
    .X(_0919_));
 sky130_fd_sc_hd__and2_1 _6560_ (.A(net858),
    .B(net171),
    .X(_0920_));
 sky130_fd_sc_hd__and2_1 _6561_ (.A(net611),
    .B(net171),
    .X(_0921_));
 sky130_fd_sc_hd__and2_1 _6562_ (.A(net742),
    .B(net172),
    .X(_0922_));
 sky130_fd_sc_hd__and2_1 _6563_ (.A(net837),
    .B(net172),
    .X(_0923_));
 sky130_fd_sc_hd__and2_1 _6564_ (.A(net798),
    .B(net172),
    .X(_0924_));
 sky130_fd_sc_hd__and2_1 _6565_ (.A(net565),
    .B(net171),
    .X(_0925_));
 sky130_fd_sc_hd__a31o_1 _6566_ (.A1(net2029),
    .A2(net919),
    .A3(_2032_),
    .B1(_2462_),
    .X(_3441_));
 sky130_fd_sc_hd__o21a_1 _6567_ (.A1(_2038_),
    .A2(_3441_),
    .B1(net175),
    .X(_0926_));
 sky130_fd_sc_hd__o211a_1 _6568_ (.A1(_1281_),
    .A2(_2034_),
    .B1(_2038_),
    .C1(net175),
    .X(_0927_));
 sky130_fd_sc_hd__and2_1 _6569_ (.A(net176),
    .B(_2448_),
    .X(_0928_));
 sky130_fd_sc_hd__o211a_1 _6570_ (.A1(_0068_),
    .A2(_2475_),
    .B1(_2465_),
    .C1(_2463_),
    .X(_3442_));
 sky130_fd_sc_hd__and3_1 _6571_ (.A(net176),
    .B(_2666_),
    .C(_3442_),
    .X(_0929_));
 sky130_fd_sc_hd__and3b_1 _6572_ (.A_N(net919),
    .B(net2037),
    .C(net2076),
    .X(_3443_));
 sky130_fd_sc_hd__and3_1 _6573_ (.A(_1280_),
    .B(_1281_),
    .C(_3443_),
    .X(_3444_));
 sky130_fd_sc_hd__a221o_1 _6574_ (.A1(_1282_),
    .A2(_2034_),
    .B1(_2462_),
    .B2(net919),
    .C1(_3444_),
    .X(_3445_));
 sky130_fd_sc_hd__o21a_1 _6575_ (.A1(_2506_),
    .A2(_3445_),
    .B1(net175),
    .X(_0930_));
 sky130_fd_sc_hd__nand2_2 _6576_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_3446_));
 sky130_fd_sc_hd__and3_2 _6577_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(net323),
    .X(_3447_));
 sky130_fd_sc_hd__inv_2 _6578_ (.A(net275),
    .Y(_3448_));
 sky130_fd_sc_hd__nor2_1 _6579_ (.A(net465),
    .B(net275),
    .Y(_3449_));
 sky130_fd_sc_hd__or2_1 _6580_ (.A(net465),
    .B(net275),
    .X(_3450_));
 sky130_fd_sc_hd__a22o_1 _6581_ (.A1(net298),
    .A2(net275),
    .B1(net229),
    .B2(net1169),
    .X(_0931_));
 sky130_fd_sc_hd__a22o_1 _6582_ (.A1(net299),
    .A2(net275),
    .B1(net229),
    .B2(net1351),
    .X(_0932_));
 sky130_fd_sc_hd__o22a_1 _6583_ (.A1(net353),
    .A2(_3448_),
    .B1(_3450_),
    .B2(net1047),
    .X(_0933_));
 sky130_fd_sc_hd__o22a_1 _6584_ (.A1(net355),
    .A2(_3448_),
    .B1(_3450_),
    .B2(net1032),
    .X(_0934_));
 sky130_fd_sc_hd__a22o_1 _6585_ (.A1(net356),
    .A2(net275),
    .B1(net229),
    .B2(net1475),
    .X(_0935_));
 sky130_fd_sc_hd__a22o_1 _6586_ (.A1(net354),
    .A2(net275),
    .B1(net229),
    .B2(net1427),
    .X(_0936_));
 sky130_fd_sc_hd__a22o_1 _6587_ (.A1(net352),
    .A2(net276),
    .B1(net228),
    .B2(net1325),
    .X(_0937_));
 sky130_fd_sc_hd__a22o_1 _6588_ (.A1(net351),
    .A2(net275),
    .B1(net228),
    .B2(net1419),
    .X(_0938_));
 sky130_fd_sc_hd__a22o_1 _6589_ (.A1(net358),
    .A2(net275),
    .B1(net229),
    .B2(net1379),
    .X(_0939_));
 sky130_fd_sc_hd__a22o_1 _6590_ (.A1(net359),
    .A2(net275),
    .B1(net229),
    .B2(net1035),
    .X(_0940_));
 sky130_fd_sc_hd__a22o_1 _6591_ (.A1(net357),
    .A2(net276),
    .B1(net228),
    .B2(net1725),
    .X(_0941_));
 sky130_fd_sc_hd__a22o_1 _6592_ (.A1(net361),
    .A2(net276),
    .B1(net228),
    .B2(net1236),
    .X(_0942_));
 sky130_fd_sc_hd__a22o_1 _6593_ (.A1(_1349_),
    .A2(net275),
    .B1(net229),
    .B2(net1678),
    .X(_0943_));
 sky130_fd_sc_hd__a22o_1 _6594_ (.A1(net360),
    .A2(net276),
    .B1(net228),
    .B2(net1262),
    .X(_0944_));
 sky130_fd_sc_hd__a22o_1 _6595_ (.A1(net350),
    .A2(net275),
    .B1(net229),
    .B2(net1563),
    .X(_0945_));
 sky130_fd_sc_hd__a22o_1 _6596_ (.A1(net349),
    .A2(_3447_),
    .B1(net229),
    .B2(net1244),
    .X(_0946_));
 sky130_fd_sc_hd__a22o_1 _6597_ (.A1(net345),
    .A2(net275),
    .B1(net229),
    .B2(net1742),
    .X(_0947_));
 sky130_fd_sc_hd__a22o_1 _6598_ (.A1(net344),
    .A2(net275),
    .B1(net229),
    .B2(net1828),
    .X(_0948_));
 sky130_fd_sc_hd__a22o_1 _6599_ (.A1(net341),
    .A2(net275),
    .B1(net229),
    .B2(net1660),
    .X(_0949_));
 sky130_fd_sc_hd__a22o_1 _6600_ (.A1(net343),
    .A2(net276),
    .B1(net228),
    .B2(net1801),
    .X(_0950_));
 sky130_fd_sc_hd__a22o_1 _6601_ (.A1(net342),
    .A2(net276),
    .B1(net228),
    .B2(net1053),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _6602_ (.A1(net346),
    .A2(net276),
    .B1(net228),
    .B2(net1662),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _6603_ (.A1(net348),
    .A2(net275),
    .B1(net229),
    .B2(net1453),
    .X(_0953_));
 sky130_fd_sc_hd__a22o_1 _6604_ (.A1(net347),
    .A2(net276),
    .B1(net228),
    .B2(net1141),
    .X(_0954_));
 sky130_fd_sc_hd__a22o_1 _6605_ (.A1(net334),
    .A2(_3447_),
    .B1(net229),
    .B2(net1617),
    .X(_0955_));
 sky130_fd_sc_hd__a22o_1 _6606_ (.A1(net337),
    .A2(net276),
    .B1(net228),
    .B2(net1153),
    .X(_0956_));
 sky130_fd_sc_hd__a22o_1 _6607_ (.A1(net338),
    .A2(net276),
    .B1(net228),
    .B2(net1479),
    .X(_0957_));
 sky130_fd_sc_hd__a22o_1 _6608_ (.A1(net336),
    .A2(net276),
    .B1(net228),
    .B2(net1545),
    .X(_0958_));
 sky130_fd_sc_hd__a22o_1 _6609_ (.A1(net333),
    .A2(net276),
    .B1(net228),
    .B2(net1511),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _6610_ (.A1(net339),
    .A2(net276),
    .B1(net228),
    .B2(net1639),
    .X(_0960_));
 sky130_fd_sc_hd__a22o_1 _6611_ (.A1(net340),
    .A2(net276),
    .B1(net228),
    .B2(net1886),
    .X(_0961_));
 sky130_fd_sc_hd__a22o_1 _6612_ (.A1(net335),
    .A2(net276),
    .B1(net228),
    .B2(net1425),
    .X(_0962_));
 sky130_fd_sc_hd__and3_2 _6613_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2620_),
    .X(_3451_));
 sky130_fd_sc_hd__nand3_2 _6614_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2620_),
    .Y(_3452_));
 sky130_fd_sc_hd__nor2_2 _6615_ (.A(net465),
    .B(net309),
    .Y(_3453_));
 sky130_fd_sc_hd__nand2_1 _6616_ (.A(net454),
    .B(_3452_),
    .Y(_3454_));
 sky130_fd_sc_hd__o22a_1 _6617_ (.A1(net298),
    .A2(_3452_),
    .B1(_3454_),
    .B2(net911),
    .X(_0963_));
 sky130_fd_sc_hd__o22a_1 _6618_ (.A1(net299),
    .A2(_3452_),
    .B1(_3454_),
    .B2(net939),
    .X(_0964_));
 sky130_fd_sc_hd__o22a_1 _6619_ (.A1(net353),
    .A2(_3452_),
    .B1(_3454_),
    .B2(net852),
    .X(_0965_));
 sky130_fd_sc_hd__o22a_1 _6620_ (.A1(net355),
    .A2(_3452_),
    .B1(_3454_),
    .B2(net935),
    .X(_0966_));
 sky130_fd_sc_hd__a22o_1 _6621_ (.A1(net356),
    .A2(net309),
    .B1(net274),
    .B2(net1688),
    .X(_0967_));
 sky130_fd_sc_hd__a22o_1 _6622_ (.A1(net354),
    .A2(net309),
    .B1(net274),
    .B2(net1381),
    .X(_0968_));
 sky130_fd_sc_hd__a22o_1 _6623_ (.A1(net352),
    .A2(net308),
    .B1(net273),
    .B2(net1615),
    .X(_0969_));
 sky130_fd_sc_hd__a22o_1 _6624_ (.A1(net351),
    .A2(net309),
    .B1(net274),
    .B2(net1723),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _6625_ (.A1(net358),
    .A2(net308),
    .B1(net273),
    .B2(net1212),
    .X(_0971_));
 sky130_fd_sc_hd__a22o_1 _6626_ (.A1(net359),
    .A2(net309),
    .B1(net274),
    .B2(net1268),
    .X(_0972_));
 sky130_fd_sc_hd__a22o_1 _6627_ (.A1(net357),
    .A2(net308),
    .B1(net273),
    .B2(net1601),
    .X(_0973_));
 sky130_fd_sc_hd__a22o_1 _6628_ (.A1(net361),
    .A2(net308),
    .B1(net273),
    .B2(net1523),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _6629_ (.A1(_1349_),
    .A2(net309),
    .B1(net274),
    .B2(net1489),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _6630_ (.A1(net360),
    .A2(net308),
    .B1(net273),
    .B2(net1059),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _6631_ (.A1(net350),
    .A2(net309),
    .B1(net274),
    .B2(net1198),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _6632_ (.A1(_1508_),
    .A2(net309),
    .B1(net274),
    .B2(net991),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _6633_ (.A1(net345),
    .A2(net309),
    .B1(net274),
    .B2(net1421),
    .X(_0979_));
 sky130_fd_sc_hd__a22o_1 _6634_ (.A1(net344),
    .A2(net309),
    .B1(net274),
    .B2(net1171),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _6635_ (.A1(net341),
    .A2(net309),
    .B1(net274),
    .B2(net1690),
    .X(_0981_));
 sky130_fd_sc_hd__a22o_1 _6636_ (.A1(net343),
    .A2(net308),
    .B1(net273),
    .B2(net1633),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _6637_ (.A1(net342),
    .A2(net308),
    .B1(net273),
    .B2(net1581),
    .X(_0983_));
 sky130_fd_sc_hd__a22o_1 _6638_ (.A1(net346),
    .A2(net308),
    .B1(net273),
    .B2(net1345),
    .X(_0984_));
 sky130_fd_sc_hd__a22o_1 _6639_ (.A1(net348),
    .A2(net309),
    .B1(net274),
    .B2(net1656),
    .X(_0985_));
 sky130_fd_sc_hd__a22o_1 _6640_ (.A1(net347),
    .A2(net308),
    .B1(net273),
    .B2(net1292),
    .X(_0986_));
 sky130_fd_sc_hd__a22o_1 _6641_ (.A1(net334),
    .A2(net309),
    .B1(net274),
    .B2(net1175),
    .X(_0987_));
 sky130_fd_sc_hd__a22o_1 _6642_ (.A1(net337),
    .A2(net308),
    .B1(net273),
    .B2(net1276),
    .X(_0988_));
 sky130_fd_sc_hd__a22o_1 _6643_ (.A1(net338),
    .A2(net308),
    .B1(net273),
    .B2(net1286),
    .X(_0989_));
 sky130_fd_sc_hd__a22o_1 _6644_ (.A1(net336),
    .A2(net308),
    .B1(net273),
    .B2(net1206),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_1 _6645_ (.A1(net333),
    .A2(net308),
    .B1(net273),
    .B2(net1539),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _6646_ (.A1(net339),
    .A2(net308),
    .B1(net273),
    .B2(net1415),
    .X(_0992_));
 sky130_fd_sc_hd__a22o_1 _6647_ (.A1(net340),
    .A2(net308),
    .B1(net273),
    .B2(net1531),
    .X(_0993_));
 sky130_fd_sc_hd__a22o_1 _6648_ (.A1(net335),
    .A2(net308),
    .B1(net273),
    .B2(net1389),
    .X(_0994_));
 sky130_fd_sc_hd__nor2_4 _6649_ (.A(_2544_),
    .B(_3446_),
    .Y(_3455_));
 sky130_fd_sc_hd__or2_2 _6650_ (.A(_2544_),
    .B(_3446_),
    .X(_3456_));
 sky130_fd_sc_hd__nor2_2 _6651_ (.A(net464),
    .B(net272),
    .Y(_3457_));
 sky130_fd_sc_hd__nand2_1 _6652_ (.A(net454),
    .B(_3456_),
    .Y(_3458_));
 sky130_fd_sc_hd__a22o_1 _6653_ (.A1(net298),
    .A2(net272),
    .B1(net227),
    .B2(net1093),
    .X(_0995_));
 sky130_fd_sc_hd__o22a_1 _6654_ (.A1(net299),
    .A2(_3456_),
    .B1(_3458_),
    .B2(net959),
    .X(_0996_));
 sky130_fd_sc_hd__o22a_1 _6655_ (.A1(net353),
    .A2(_3456_),
    .B1(_3458_),
    .B2(net901),
    .X(_0997_));
 sky130_fd_sc_hd__o22a_1 _6656_ (.A1(net355),
    .A2(_3456_),
    .B1(_3458_),
    .B2(net947),
    .X(_0998_));
 sky130_fd_sc_hd__a22o_1 _6657_ (.A1(net356),
    .A2(net272),
    .B1(net227),
    .B2(net1327),
    .X(_0999_));
 sky130_fd_sc_hd__a22o_1 _6658_ (.A1(net354),
    .A2(net272),
    .B1(net227),
    .B2(net1795),
    .X(_1000_));
 sky130_fd_sc_hd__a22o_1 _6659_ (.A1(net352),
    .A2(net271),
    .B1(net226),
    .B2(net1585),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _6660_ (.A1(net351),
    .A2(net271),
    .B1(net227),
    .B2(net1367),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _6661_ (.A1(net358),
    .A2(net272),
    .B1(net226),
    .B2(net1123),
    .X(_1003_));
 sky130_fd_sc_hd__a22o_1 _6662_ (.A1(net359),
    .A2(net272),
    .B1(net227),
    .B2(net1248),
    .X(_1004_));
 sky130_fd_sc_hd__a22o_1 _6663_ (.A1(net357),
    .A2(net271),
    .B1(net226),
    .B2(net1437),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _6664_ (.A1(net361),
    .A2(net271),
    .B1(net226),
    .B2(net1635),
    .X(_1006_));
 sky130_fd_sc_hd__a22o_1 _6665_ (.A1(_1349_),
    .A2(net272),
    .B1(net227),
    .B2(net1391),
    .X(_1007_));
 sky130_fd_sc_hd__a22o_1 _6666_ (.A1(net360),
    .A2(net271),
    .B1(net226),
    .B2(net1625),
    .X(_1008_));
 sky130_fd_sc_hd__a22o_1 _6667_ (.A1(net350),
    .A2(net272),
    .B1(net227),
    .B2(net1252),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _6668_ (.A1(net349),
    .A2(net272),
    .B1(net227),
    .B2(net1228),
    .X(_1010_));
 sky130_fd_sc_hd__a22o_1 _6669_ (.A1(net345),
    .A2(net272),
    .B1(net227),
    .B2(net1469),
    .X(_1011_));
 sky130_fd_sc_hd__a22o_1 _6670_ (.A1(net344),
    .A2(net272),
    .B1(net227),
    .B2(net1008),
    .X(_1012_));
 sky130_fd_sc_hd__a22o_1 _6671_ (.A1(net341),
    .A2(net272),
    .B1(net227),
    .B2(net1481),
    .X(_1013_));
 sky130_fd_sc_hd__a22o_1 _6672_ (.A1(net343),
    .A2(net271),
    .B1(net226),
    .B2(net1463),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _6673_ (.A1(net342),
    .A2(net271),
    .B1(net226),
    .B2(net1455),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_1 _6674_ (.A1(net346),
    .A2(net271),
    .B1(net226),
    .B2(net1781),
    .X(_1016_));
 sky130_fd_sc_hd__a22o_1 _6675_ (.A1(net348),
    .A2(net272),
    .B1(net227),
    .B2(net1735),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _6676_ (.A1(net347),
    .A2(net271),
    .B1(net226),
    .B2(net1234),
    .X(_1018_));
 sky130_fd_sc_hd__a22o_1 _6677_ (.A1(net334),
    .A2(net272),
    .B1(net227),
    .B2(net1694),
    .X(_1019_));
 sky130_fd_sc_hd__a22o_1 _6678_ (.A1(net337),
    .A2(net271),
    .B1(net226),
    .B2(net1501),
    .X(_1020_));
 sky130_fd_sc_hd__a22o_1 _6679_ (.A1(net338),
    .A2(net271),
    .B1(net226),
    .B2(net1429),
    .X(_1021_));
 sky130_fd_sc_hd__a22o_1 _6680_ (.A1(net336),
    .A2(net271),
    .B1(net226),
    .B2(net1242),
    .X(_1022_));
 sky130_fd_sc_hd__a22o_1 _6681_ (.A1(net333),
    .A2(net271),
    .B1(net226),
    .B2(net1573),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _6682_ (.A1(net339),
    .A2(net271),
    .B1(net226),
    .B2(net1449),
    .X(_1024_));
 sky130_fd_sc_hd__a22o_1 _6683_ (.A1(net340),
    .A2(net271),
    .B1(net226),
    .B2(net1264),
    .X(_1025_));
 sky130_fd_sc_hd__a22o_1 _6684_ (.A1(_1632_),
    .A2(net271),
    .B1(net226),
    .B2(net1485),
    .X(_1026_));
 sky130_fd_sc_hd__nor2_1 _6685_ (.A(_2509_),
    .B(_2626_),
    .Y(_3459_));
 sky130_fd_sc_hd__or2_1 _6686_ (.A(_2509_),
    .B(_2626_),
    .X(_3460_));
 sky130_fd_sc_hd__nor2_1 _6687_ (.A(net465),
    .B(net270),
    .Y(_3461_));
 sky130_fd_sc_hd__nand2_1 _6688_ (.A(net447),
    .B(_3460_),
    .Y(_3462_));
 sky130_fd_sc_hd__o22a_1 _6689_ (.A1(net298),
    .A2(_3460_),
    .B1(_3462_),
    .B2(net893),
    .X(_1027_));
 sky130_fd_sc_hd__a22o_1 _6690_ (.A1(net299),
    .A2(net270),
    .B1(net225),
    .B2(net1699),
    .X(_1028_));
 sky130_fd_sc_hd__o22a_1 _6691_ (.A1(net353),
    .A2(_3460_),
    .B1(_3462_),
    .B2(net925),
    .X(_1029_));
 sky130_fd_sc_hd__a22o_1 _6692_ (.A1(net355),
    .A2(net270),
    .B1(net225),
    .B2(net1565),
    .X(_1030_));
 sky130_fd_sc_hd__a22o_1 _6693_ (.A1(net356),
    .A2(net270),
    .B1(net225),
    .B2(net1091),
    .X(_1031_));
 sky130_fd_sc_hd__a22o_1 _6694_ (.A1(net354),
    .A2(net270),
    .B1(net225),
    .B2(net1069),
    .X(_1032_));
 sky130_fd_sc_hd__a22o_1 _6695_ (.A1(net352),
    .A2(net269),
    .B1(net224),
    .B2(net1567),
    .X(_1033_));
 sky130_fd_sc_hd__a22o_1 _6696_ (.A1(net351),
    .A2(net269),
    .B1(net224),
    .B2(net1129),
    .X(_1034_));
 sky130_fd_sc_hd__a22o_1 _6697_ (.A1(net358),
    .A2(net269),
    .B1(net224),
    .B2(net1411),
    .X(_1035_));
 sky130_fd_sc_hd__a22o_1 _6698_ (.A1(net359),
    .A2(net270),
    .B1(net225),
    .B2(net965),
    .X(_1036_));
 sky130_fd_sc_hd__a22o_1 _6699_ (.A1(net357),
    .A2(net269),
    .B1(net224),
    .B2(net1173),
    .X(_1037_));
 sky130_fd_sc_hd__a22o_1 _6700_ (.A1(net361),
    .A2(net269),
    .B1(net224),
    .B2(net1547),
    .X(_1038_));
 sky130_fd_sc_hd__a22o_1 _6701_ (.A1(_1349_),
    .A2(net270),
    .B1(net225),
    .B2(net1022),
    .X(_1039_));
 sky130_fd_sc_hd__a22o_1 _6702_ (.A1(net360),
    .A2(net269),
    .B1(net224),
    .B2(net1322),
    .X(_1040_));
 sky130_fd_sc_hd__a22o_1 _6703_ (.A1(net350),
    .A2(net270),
    .B1(net225),
    .B2(net1111),
    .X(_1041_));
 sky130_fd_sc_hd__a22o_1 _6704_ (.A1(net349),
    .A2(net270),
    .B1(net225),
    .B2(net1457),
    .X(_1042_));
 sky130_fd_sc_hd__a22o_1 _6705_ (.A1(net345),
    .A2(net270),
    .B1(net225),
    .B2(net1159),
    .X(_1043_));
 sky130_fd_sc_hd__a22o_1 _6706_ (.A1(net344),
    .A2(net270),
    .B1(net225),
    .B2(net1294),
    .X(_1044_));
 sky130_fd_sc_hd__a22o_1 _6707_ (.A1(net341),
    .A2(net270),
    .B1(net225),
    .B2(net1593),
    .X(_1045_));
 sky130_fd_sc_hd__a22o_1 _6708_ (.A1(net343),
    .A2(net269),
    .B1(net224),
    .B2(net1185),
    .X(_1046_));
 sky130_fd_sc_hd__a22o_1 _6709_ (.A1(net342),
    .A2(net269),
    .B1(net224),
    .B2(net1065),
    .X(_1047_));
 sky130_fd_sc_hd__a22o_1 _6710_ (.A1(net346),
    .A2(net269),
    .B1(net224),
    .B2(net1179),
    .X(_1048_));
 sky130_fd_sc_hd__a22o_1 _6711_ (.A1(net348),
    .A2(net270),
    .B1(net225),
    .B2(net1081),
    .X(_1049_));
 sky130_fd_sc_hd__a22o_1 _6712_ (.A1(net347),
    .A2(net269),
    .B1(net224),
    .B2(net1099),
    .X(_1050_));
 sky130_fd_sc_hd__a22o_1 _6713_ (.A1(net334),
    .A2(net270),
    .B1(net225),
    .B2(net1533),
    .X(_1051_));
 sky130_fd_sc_hd__a22o_1 _6714_ (.A1(net337),
    .A2(net269),
    .B1(net224),
    .B2(net1709),
    .X(_1052_));
 sky130_fd_sc_hd__a22o_1 _6715_ (.A1(net338),
    .A2(net269),
    .B1(net224),
    .B2(net1061),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_1 _6716_ (.A1(net336),
    .A2(net270),
    .B1(net225),
    .B2(net1020),
    .X(_1054_));
 sky130_fd_sc_hd__a22o_1 _6717_ (.A1(net333),
    .A2(net269),
    .B1(net224),
    .B2(net1214),
    .X(_1055_));
 sky130_fd_sc_hd__a22o_1 _6718_ (.A1(net339),
    .A2(net269),
    .B1(net224),
    .B2(net945),
    .X(_1056_));
 sky130_fd_sc_hd__a22o_1 _6719_ (.A1(net340),
    .A2(net269),
    .B1(net224),
    .B2(net997),
    .X(_1057_));
 sky130_fd_sc_hd__a22o_1 _6720_ (.A1(net335),
    .A2(net269),
    .B1(net224),
    .B2(net1571),
    .X(_1058_));
 sky130_fd_sc_hd__and2_1 _6721_ (.A(net454),
    .B(net1079),
    .X(_1059_));
 sky130_fd_sc_hd__and2_1 _6722_ (.A(net447),
    .B(net1005),
    .X(_1060_));
 sky130_fd_sc_hd__and2_1 _6723_ (.A(net447),
    .B(net1587),
    .X(_1061_));
 sky130_fd_sc_hd__and2_1 _6724_ (.A(net455),
    .B(net1431),
    .X(_1062_));
 sky130_fd_sc_hd__and2_1 _6725_ (.A(net455),
    .B(net1497),
    .X(_1063_));
 sky130_fd_sc_hd__and2_1 _6726_ (.A(net452),
    .B(net1525),
    .X(_1064_));
 sky130_fd_sc_hd__and2_1 _6727_ (.A(net439),
    .B(net1290),
    .X(_1065_));
 sky130_fd_sc_hd__and2_1 _6728_ (.A(net445),
    .B(net1192),
    .X(_1066_));
 sky130_fd_sc_hd__and2_1 _6729_ (.A(net446),
    .B(net1529),
    .X(_1067_));
 sky130_fd_sc_hd__and2_1 _6730_ (.A(net456),
    .B(net1553),
    .X(_1068_));
 sky130_fd_sc_hd__and2_1 _6731_ (.A(net439),
    .B(net1637),
    .X(_1069_));
 sky130_fd_sc_hd__and2_1 _6732_ (.A(net430),
    .B(net1549),
    .X(_1070_));
 sky130_fd_sc_hd__and2_1 _6733_ (.A(net452),
    .B(net1527),
    .X(_1071_));
 sky130_fd_sc_hd__and2_1 _6734_ (.A(net439),
    .B(net1238),
    .X(_1072_));
 sky130_fd_sc_hd__and2_1 _6735_ (.A(net451),
    .B(net1599),
    .X(_1073_));
 sky130_fd_sc_hd__and2_1 _6736_ (.A(net442),
    .B(net1151),
    .X(_1074_));
 sky130_fd_sc_hd__and2_1 _6737_ (.A(net445),
    .B(net1024),
    .X(_1075_));
 sky130_fd_sc_hd__and2_1 _6738_ (.A(net448),
    .B(net1621),
    .X(_1076_));
 sky130_fd_sc_hd__and2_1 _6739_ (.A(net455),
    .B(net1748),
    .X(_1077_));
 sky130_fd_sc_hd__and2_1 _6740_ (.A(net438),
    .B(net1793),
    .X(_1078_));
 sky130_fd_sc_hd__and2_1 _6741_ (.A(net436),
    .B(net1401),
    .X(_1079_));
 sky130_fd_sc_hd__and2_1 _6742_ (.A(net437),
    .B(net1676),
    .X(_1080_));
 sky130_fd_sc_hd__and2_1 _6743_ (.A(net445),
    .B(net1439),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _6744_ (.A(net434),
    .B(net1077),
    .X(_1082_));
 sky130_fd_sc_hd__and2_1 _6745_ (.A(net455),
    .B(net1649),
    .X(_1083_));
 sky130_fd_sc_hd__and2_1 _6746_ (.A(net433),
    .B(net1254),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _6747_ (.A(net434),
    .B(net1073),
    .X(_1085_));
 sky130_fd_sc_hd__and2_1 _6748_ (.A(net438),
    .B(net1399),
    .X(_1086_));
 sky130_fd_sc_hd__and2_1 _6749_ (.A(net430),
    .B(net1026),
    .X(_1087_));
 sky130_fd_sc_hd__and2_1 _6750_ (.A(net433),
    .B(net1385),
    .X(_1088_));
 sky130_fd_sc_hd__and2_1 _6751_ (.A(net436),
    .B(net1447),
    .X(_1089_));
 sky130_fd_sc_hd__and2_1 _6752_ (.A(net434),
    .B(net1721),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_1 _6753_ (.A(_2544_),
    .B(_2626_),
    .Y(_3463_));
 sky130_fd_sc_hd__or2_2 _6754_ (.A(_2544_),
    .B(_2626_),
    .X(_3464_));
 sky130_fd_sc_hd__nor2_1 _6755_ (.A(net465),
    .B(net268),
    .Y(_3465_));
 sky130_fd_sc_hd__nand2_1 _6756_ (.A(net447),
    .B(_3464_),
    .Y(_3466_));
 sky130_fd_sc_hd__a22o_1 _6757_ (.A1(net298),
    .A2(net268),
    .B1(net223),
    .B2(net1310),
    .X(_1091_));
 sky130_fd_sc_hd__o22a_1 _6758_ (.A1(_1440_),
    .A2(_3464_),
    .B1(_3466_),
    .B2(net995),
    .X(_1092_));
 sky130_fd_sc_hd__o22a_1 _6759_ (.A1(net353),
    .A2(_3464_),
    .B1(_3466_),
    .B2(net871),
    .X(_1093_));
 sky130_fd_sc_hd__a22o_1 _6760_ (.A1(net355),
    .A2(net268),
    .B1(net223),
    .B2(net987),
    .X(_1094_));
 sky130_fd_sc_hd__a22o_1 _6761_ (.A1(_1420_),
    .A2(net268),
    .B1(net223),
    .B2(net1256),
    .X(_1095_));
 sky130_fd_sc_hd__a22o_1 _6762_ (.A1(_1453_),
    .A2(net268),
    .B1(net223),
    .B2(net1139),
    .X(_1096_));
 sky130_fd_sc_hd__a22o_1 _6763_ (.A1(net352),
    .A2(net267),
    .B1(net222),
    .B2(net1623),
    .X(_1097_));
 sky130_fd_sc_hd__a22o_1 _6764_ (.A1(net351),
    .A2(net268),
    .B1(net223),
    .B2(net1230),
    .X(_1098_));
 sky130_fd_sc_hd__a22o_1 _6765_ (.A1(net358),
    .A2(net267),
    .B1(net222),
    .B2(net1202),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_1 _6766_ (.A1(net359),
    .A2(net268),
    .B1(net223),
    .B2(net1095),
    .X(_1100_));
 sky130_fd_sc_hd__a22o_1 _6767_ (.A1(net357),
    .A2(net267),
    .B1(net222),
    .B2(net1204),
    .X(_1101_));
 sky130_fd_sc_hd__a22o_1 _6768_ (.A1(net361),
    .A2(net267),
    .B1(net222),
    .B2(net1147),
    .X(_1102_));
 sky130_fd_sc_hd__a22o_1 _6769_ (.A1(_1349_),
    .A2(net268),
    .B1(net223),
    .B2(net1561),
    .X(_1103_));
 sky130_fd_sc_hd__a22o_1 _6770_ (.A1(net360),
    .A2(net267),
    .B1(net222),
    .B2(net1196),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _6771_ (.A1(net350),
    .A2(net268),
    .B1(net223),
    .B2(net1067),
    .X(_1105_));
 sky130_fd_sc_hd__a22o_1 _6772_ (.A1(net349),
    .A2(net268),
    .B1(net223),
    .B2(net1274),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _6773_ (.A1(net345),
    .A2(net268),
    .B1(net223),
    .B2(net1012),
    .X(_1107_));
 sky130_fd_sc_hd__a22o_1 _6774_ (.A1(_1554_),
    .A2(net268),
    .B1(net223),
    .B2(net1609),
    .X(_1108_));
 sky130_fd_sc_hd__a22o_1 _6775_ (.A1(_1579_),
    .A2(net268),
    .B1(net223),
    .B2(net1320),
    .X(_1109_));
 sky130_fd_sc_hd__a22o_1 _6776_ (.A1(net343),
    .A2(net267),
    .B1(net222),
    .B2(net1641),
    .X(_1110_));
 sky130_fd_sc_hd__a22o_1 _6777_ (.A1(_1569_),
    .A2(net267),
    .B1(net222),
    .B2(net1157),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _6778_ (.A1(net346),
    .A2(net267),
    .B1(net222),
    .B2(net1210),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _6779_ (.A1(net348),
    .A2(net268),
    .B1(net223),
    .B2(net1075),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_1 _6780_ (.A1(net347),
    .A2(net267),
    .B1(net222),
    .B2(net1551),
    .X(_1114_));
 sky130_fd_sc_hd__a22o_1 _6781_ (.A1(net334),
    .A2(net268),
    .B1(net223),
    .B2(net1339),
    .X(_1115_));
 sky130_fd_sc_hd__a22o_1 _6782_ (.A1(net337),
    .A2(net267),
    .B1(net222),
    .B2(net1702),
    .X(_1116_));
 sky130_fd_sc_hd__a22o_1 _6783_ (.A1(net338),
    .A2(net267),
    .B1(net222),
    .B2(net1589),
    .X(_1117_));
 sky130_fd_sc_hd__a22o_1 _6784_ (.A1(net336),
    .A2(net267),
    .B1(net222),
    .B2(net1003),
    .X(_1118_));
 sky130_fd_sc_hd__a22o_1 _6785_ (.A1(net333),
    .A2(net267),
    .B1(net222),
    .B2(net1341),
    .X(_1119_));
 sky130_fd_sc_hd__a22o_1 _6786_ (.A1(net339),
    .A2(net267),
    .B1(net222),
    .B2(net1109),
    .X(_1120_));
 sky130_fd_sc_hd__a22o_1 _6787_ (.A1(net340),
    .A2(net267),
    .B1(net222),
    .B2(net1433),
    .X(_1121_));
 sky130_fd_sc_hd__a22o_1 _6788_ (.A1(net335),
    .A2(net267),
    .B1(net222),
    .B2(net1107),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_2 _6789_ (.A(_2509_),
    .B(_3446_),
    .Y(_3467_));
 sky130_fd_sc_hd__or2_1 _6790_ (.A(_2509_),
    .B(_3446_),
    .X(_3468_));
 sky130_fd_sc_hd__nor2_1 _6791_ (.A(net464),
    .B(net307),
    .Y(_3469_));
 sky130_fd_sc_hd__nand2_1 _6792_ (.A(net454),
    .B(_3468_),
    .Y(_3470_));
 sky130_fd_sc_hd__o22a_1 _6793_ (.A1(_1472_),
    .A2(_3468_),
    .B1(_3470_),
    .B2(net917),
    .X(_1123_));
 sky130_fd_sc_hd__a22o_1 _6794_ (.A1(net299),
    .A2(net307),
    .B1(net266),
    .B2(net1284),
    .X(_1124_));
 sky130_fd_sc_hd__o22a_1 _6795_ (.A1(net353),
    .A2(_3468_),
    .B1(_3470_),
    .B2(net1423),
    .X(_1125_));
 sky130_fd_sc_hd__o22a_1 _6796_ (.A1(_1430_),
    .A2(_3468_),
    .B1(_3470_),
    .B2(net867),
    .X(_1126_));
 sky130_fd_sc_hd__a22o_1 _6797_ (.A1(net356),
    .A2(net307),
    .B1(net266),
    .B2(net1733),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _6798_ (.A1(net354),
    .A2(net307),
    .B1(net266),
    .B2(net1103),
    .X(_1128_));
 sky130_fd_sc_hd__a22o_1 _6799_ (.A1(net352),
    .A2(net306),
    .B1(net265),
    .B2(net1119),
    .X(_1129_));
 sky130_fd_sc_hd__a22o_1 _6800_ (.A1(net351),
    .A2(net307),
    .B1(net266),
    .B2(net1445),
    .X(_1130_));
 sky130_fd_sc_hd__a22o_1 _6801_ (.A1(_1402_),
    .A2(net306),
    .B1(net265),
    .B2(net1495),
    .X(_1131_));
 sky130_fd_sc_hd__a22o_1 _6802_ (.A1(_1392_),
    .A2(net307),
    .B1(net266),
    .B2(net1045),
    .X(_1132_));
 sky130_fd_sc_hd__a22o_1 _6803_ (.A1(_1412_),
    .A2(net306),
    .B1(net265),
    .B2(net1707),
    .X(_1133_));
 sky130_fd_sc_hd__a22o_1 _6804_ (.A1(net361),
    .A2(net306),
    .B1(net265),
    .B2(net927),
    .X(_1134_));
 sky130_fd_sc_hd__a22o_1 _6805_ (.A1(_1349_),
    .A2(net307),
    .B1(net266),
    .B2(net1866),
    .X(_1135_));
 sky130_fd_sc_hd__a22o_1 _6806_ (.A1(_1384_),
    .A2(net306),
    .B1(net265),
    .B2(net1403),
    .X(_1136_));
 sky130_fd_sc_hd__a22o_1 _6807_ (.A1(_1501_),
    .A2(net307),
    .B1(net266),
    .B2(net1559),
    .X(_1137_));
 sky130_fd_sc_hd__a22o_1 _6808_ (.A1(net349),
    .A2(net307),
    .B1(net266),
    .B2(net1030),
    .X(_1138_));
 sky130_fd_sc_hd__a22o_1 _6809_ (.A1(_1545_),
    .A2(net307),
    .B1(net266),
    .B2(net1377),
    .X(_1139_));
 sky130_fd_sc_hd__a22o_1 _6810_ (.A1(net344),
    .A2(net307),
    .B1(net266),
    .B2(net1597),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _6811_ (.A1(net341),
    .A2(net307),
    .B1(net266),
    .B2(net1712),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _6812_ (.A1(net343),
    .A2(net306),
    .B1(net265),
    .B2(net1347),
    .X(_1142_));
 sky130_fd_sc_hd__a22o_1 _6813_ (.A1(net342),
    .A2(net306),
    .B1(net265),
    .B2(net1187),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _6814_ (.A1(_1535_),
    .A2(net306),
    .B1(net265),
    .B2(net1407),
    .X(_1144_));
 sky130_fd_sc_hd__a22o_1 _6815_ (.A1(net348),
    .A2(net307),
    .B1(net266),
    .B2(net1393),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_1 _6816_ (.A1(net347),
    .A2(net306),
    .B1(net265),
    .B2(net951),
    .X(_1146_));
 sky130_fd_sc_hd__a22o_1 _6817_ (.A1(net334),
    .A2(net307),
    .B1(net266),
    .B2(net1658),
    .X(_1147_));
 sky130_fd_sc_hd__a22o_1 _6818_ (.A1(_1613_),
    .A2(net306),
    .B1(net265),
    .B2(net1232),
    .X(_1148_));
 sky130_fd_sc_hd__a22o_1 _6819_ (.A1(_1605_),
    .A2(net306),
    .B1(net265),
    .B2(net1016),
    .X(_1149_));
 sky130_fd_sc_hd__a22o_1 _6820_ (.A1(_1622_),
    .A2(net306),
    .B1(net265),
    .B2(net1607),
    .X(_1150_));
 sky130_fd_sc_hd__a22o_1 _6821_ (.A1(net333),
    .A2(net306),
    .B1(net265),
    .B2(net1503),
    .X(_1151_));
 sky130_fd_sc_hd__a22o_1 _6822_ (.A1(_1596_),
    .A2(net306),
    .B1(net265),
    .B2(net1441),
    .X(_1152_));
 sky130_fd_sc_hd__a22o_1 _6823_ (.A1(_1588_),
    .A2(net306),
    .B1(net265),
    .B2(net1105),
    .X(_1153_));
 sky130_fd_sc_hd__a22o_1 _6824_ (.A1(net335),
    .A2(net306),
    .B1(net265),
    .B2(net1361),
    .X(_1154_));
 sky130_fd_sc_hd__and3_1 _6825_ (.A(_1301_),
    .B(net435),
    .C(_1707_),
    .X(_3471_));
 sky130_fd_sc_hd__or2_1 _6826_ (.A(net822),
    .B(net250),
    .X(_3472_));
 sky130_fd_sc_hd__o211a_1 _6827_ (.A1(net976),
    .A2(net261),
    .B1(net170),
    .C1(_3472_),
    .X(_1155_));
 sky130_fd_sc_hd__or2_1 _6828_ (.A(net769),
    .B(net252),
    .X(_3473_));
 sky130_fd_sc_hd__o211a_1 _6829_ (.A1(net903),
    .A2(net263),
    .B1(net168),
    .C1(_3473_),
    .X(_1156_));
 sky130_fd_sc_hd__or2_1 _6830_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ),
    .B(net252),
    .X(_3474_));
 sky130_fd_sc_hd__o211a_1 _6831_ (.A1(net756),
    .A2(net263),
    .B1(net168),
    .C1(_3474_),
    .X(_1157_));
 sky130_fd_sc_hd__or2_1 _6832_ (.A(net812),
    .B(net251),
    .X(_3475_));
 sky130_fd_sc_hd__o211a_1 _6833_ (.A1(net820),
    .A2(net263),
    .B1(net168),
    .C1(_3475_),
    .X(_1158_));
 sky130_fd_sc_hd__or2_1 _6834_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ),
    .B(net250),
    .X(_3476_));
 sky130_fd_sc_hd__o211a_1 _6835_ (.A1(net787),
    .A2(net261),
    .B1(net170),
    .C1(_3476_),
    .X(_1159_));
 sky130_fd_sc_hd__or2_1 _6836_ (.A(net796),
    .B(net249),
    .X(_3477_));
 sky130_fd_sc_hd__o211a_1 _6837_ (.A1(net941),
    .A2(net259),
    .B1(net167),
    .C1(_3477_),
    .X(_1160_));
 sky130_fd_sc_hd__or2_1 _6838_ (.A(net865),
    .B(net249),
    .X(_3478_));
 sky130_fd_sc_hd__o211a_1 _6839_ (.A1(net953),
    .A2(net259),
    .B1(net167),
    .C1(_3478_),
    .X(_1161_));
 sky130_fd_sc_hd__or2_1 _6840_ (.A(net804),
    .B(net252),
    .X(_3479_));
 sky130_fd_sc_hd__o211a_1 _6841_ (.A1(net963),
    .A2(net263),
    .B1(net169),
    .C1(_3479_),
    .X(_1162_));
 sky130_fd_sc_hd__or2_1 _6842_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ),
    .B(net248),
    .X(_3480_));
 sky130_fd_sc_hd__o211a_1 _6843_ (.A1(net806),
    .A2(net258),
    .B1(net166),
    .C1(_3480_),
    .X(_1163_));
 sky130_fd_sc_hd__or2_1 _6844_ (.A(net887),
    .B(net251),
    .X(_3481_));
 sky130_fd_sc_hd__o211a_1 _6845_ (.A1(net1101),
    .A2(net262),
    .B1(net168),
    .C1(_3481_),
    .X(_1164_));
 sky130_fd_sc_hd__or2_1 _6846_ (.A(net843),
    .B(net252),
    .X(_3482_));
 sky130_fd_sc_hd__o211a_1 _6847_ (.A1(net989),
    .A2(net263),
    .B1(net168),
    .C1(_3482_),
    .X(_1165_));
 sky130_fd_sc_hd__or2_1 _6848_ (.A(net561),
    .B(net250),
    .X(_3483_));
 sky130_fd_sc_hd__o211a_1 _6849_ (.A1(net905),
    .A2(net261),
    .B1(net170),
    .C1(_3483_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_1 _6850_ (.A(net832),
    .B(net252),
    .X(_3484_));
 sky130_fd_sc_hd__o211a_1 _6851_ (.A1(net1001),
    .A2(net263),
    .B1(net169),
    .C1(_3484_),
    .X(_1167_));
 sky130_fd_sc_hd__or2_1 _6852_ (.A(net571),
    .B(net251),
    .X(_3485_));
 sky130_fd_sc_hd__o211a_1 _6853_ (.A1(net1083),
    .A2(net262),
    .B1(net168),
    .C1(_3485_),
    .X(_1168_));
 sky130_fd_sc_hd__or2_1 _6854_ (.A(net541),
    .B(net250),
    .X(_3486_));
 sky130_fd_sc_hd__o211a_1 _6855_ (.A1(net915),
    .A2(net259),
    .B1(net167),
    .C1(_3486_),
    .X(_1169_));
 sky130_fd_sc_hd__or2_1 _6856_ (.A(net791),
    .B(net250),
    .X(_3487_));
 sky130_fd_sc_hd__o211a_1 _6857_ (.A1(net937),
    .A2(net261),
    .B1(net170),
    .C1(_3487_),
    .X(_1170_));
 sky130_fd_sc_hd__or2_1 _6858_ (.A(net609),
    .B(net252),
    .X(_3488_));
 sky130_fd_sc_hd__o211a_1 _6859_ (.A1(net981),
    .A2(net263),
    .B1(net169),
    .C1(_3488_),
    .X(_1171_));
 sky130_fd_sc_hd__or2_1 _6860_ (.A(net835),
    .B(net250),
    .X(_3489_));
 sky130_fd_sc_hd__o211a_1 _6861_ (.A1(net1143),
    .A2(net261),
    .B1(net170),
    .C1(_3489_),
    .X(_1172_));
 sky130_fd_sc_hd__or2_1 _6862_ (.A(net891),
    .B(net246),
    .X(_3490_));
 sky130_fd_sc_hd__o211a_1 _6863_ (.A1(net955),
    .A2(net255),
    .B1(net164),
    .C1(_3490_),
    .X(_1173_));
 sky130_fd_sc_hd__or2_1 _6864_ (.A(net869),
    .B(net247),
    .X(_3491_));
 sky130_fd_sc_hd__o211a_1 _6865_ (.A1(net972),
    .A2(net256),
    .B1(net164),
    .C1(_3491_),
    .X(_1174_));
 sky130_fd_sc_hd__or2_1 _6866_ (.A(net845),
    .B(net244),
    .X(_3492_));
 sky130_fd_sc_hd__o211a_1 _6867_ (.A1(net943),
    .A2(net254),
    .B1(net165),
    .C1(_3492_),
    .X(_1175_));
 sky130_fd_sc_hd__or2_1 _6868_ (.A(net897),
    .B(net244),
    .X(_3493_));
 sky130_fd_sc_hd__o211a_1 _6869_ (.A1(net923),
    .A2(net254),
    .B1(net165),
    .C1(_3493_),
    .X(_1176_));
 sky130_fd_sc_hd__or2_1 _6870_ (.A(net974),
    .B(net246),
    .X(_3494_));
 sky130_fd_sc_hd__o211a_1 _6871_ (.A1(net1043),
    .A2(net256),
    .B1(net164),
    .C1(_3494_),
    .X(_1177_));
 sky130_fd_sc_hd__or2_1 _6872_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ),
    .B(net247),
    .X(_3495_));
 sky130_fd_sc_hd__o211a_1 _6873_ (.A1(net668),
    .A2(net256),
    .B1(net164),
    .C1(_3495_),
    .X(_1178_));
 sky130_fd_sc_hd__or2_1 _6874_ (.A(net883),
    .B(net247),
    .X(_3496_));
 sky130_fd_sc_hd__o211a_1 _6875_ (.A1(net1018),
    .A2(net256),
    .B1(net164),
    .C1(_3496_),
    .X(_1179_));
 sky130_fd_sc_hd__or2_1 _6876_ (.A(net644),
    .B(net245),
    .X(_3497_));
 sky130_fd_sc_hd__o211a_1 _6877_ (.A1(net929),
    .A2(net254),
    .B1(net165),
    .C1(_3497_),
    .X(_1180_));
 sky130_fd_sc_hd__or2_1 _6878_ (.A(net879),
    .B(net244),
    .X(_3498_));
 sky130_fd_sc_hd__o211a_1 _6879_ (.A1(net913),
    .A2(net254),
    .B1(net165),
    .C1(_3498_),
    .X(_1181_));
 sky130_fd_sc_hd__or2_1 _6880_ (.A(net563),
    .B(net245),
    .X(_3499_));
 sky130_fd_sc_hd__o211a_1 _6881_ (.A1(net854),
    .A2(net254),
    .B1(net165),
    .C1(_3499_),
    .X(_1182_));
 sky130_fd_sc_hd__or2_1 _6882_ (.A(net800),
    .B(net245),
    .X(_3500_));
 sky130_fd_sc_hd__o211a_1 _6883_ (.A1(net933),
    .A2(net257),
    .B1(net165),
    .C1(_3500_),
    .X(_1183_));
 sky130_fd_sc_hd__or2_1 _6884_ (.A(net818),
    .B(net248),
    .X(_3501_));
 sky130_fd_sc_hd__o211a_1 _6885_ (.A1(net899),
    .A2(net257),
    .B1(net166),
    .C1(_3501_),
    .X(_1184_));
 sky130_fd_sc_hd__or2_1 _6886_ (.A(net2076),
    .B(net245),
    .X(_3502_));
 sky130_fd_sc_hd__o211a_1 _6887_ (.A1(net21),
    .A2(net257),
    .B1(net165),
    .C1(_3502_),
    .X(_1185_));
 sky130_fd_sc_hd__or2_1 _6888_ (.A(net2037),
    .B(net249),
    .X(_3503_));
 sky130_fd_sc_hd__o211a_1 _6889_ (.A1(net24),
    .A2(net259),
    .B1(net167),
    .C1(_3503_),
    .X(_1186_));
 sky130_fd_sc_hd__mux2_1 _6890_ (.A0(net25),
    .A1(net919),
    .S(net260),
    .X(_3504_));
 sky130_fd_sc_hd__nand2b_1 _6891_ (.A_N(_3504_),
    .B(net167),
    .Y(_1187_));
 sky130_fd_sc_hd__nand2_1 _6892_ (.A(net26),
    .B(net249),
    .Y(_3505_));
 sky130_fd_sc_hd__o211ai_1 _6893_ (.A1(_1281_),
    .A2(net249),
    .B1(net167),
    .C1(_3505_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _6894_ (.A(_1280_),
    .B(net260),
    .Y(_3506_));
 sky130_fd_sc_hd__o211a_1 _6895_ (.A1(net27),
    .A2(net260),
    .B1(net167),
    .C1(_3506_),
    .X(_1189_));
 sky130_fd_sc_hd__or2_1 _6896_ (.A(net1959),
    .B(net252),
    .X(_3507_));
 sky130_fd_sc_hd__o211a_1 _6897_ (.A1(net28),
    .A2(net263),
    .B1(net168),
    .C1(_3507_),
    .X(_1190_));
 sky130_fd_sc_hd__or2_1 _6898_ (.A(net1946),
    .B(net249),
    .X(_3508_));
 sky130_fd_sc_hd__o211a_1 _6899_ (.A1(net29),
    .A2(net259),
    .B1(net167),
    .C1(_3508_),
    .X(_1191_));
 sky130_fd_sc_hd__or2_1 _6900_ (.A(net2042),
    .B(net253),
    .X(_3509_));
 sky130_fd_sc_hd__o211a_1 _6901_ (.A1(net30),
    .A2(net264),
    .B1(net169),
    .C1(_3509_),
    .X(_1192_));
 sky130_fd_sc_hd__or2_1 _6902_ (.A(net608),
    .B(net253),
    .X(_3510_));
 sky130_fd_sc_hd__o211a_1 _6903_ (.A1(net1),
    .A2(net263),
    .B1(net168),
    .C1(_3510_),
    .X(_1193_));
 sky130_fd_sc_hd__or2_1 _6904_ (.A(net2127),
    .B(net248),
    .X(_3511_));
 sky130_fd_sc_hd__o211a_1 _6905_ (.A1(net2),
    .A2(net258),
    .B1(net166),
    .C1(_3511_),
    .X(_1194_));
 sky130_fd_sc_hd__or2_1 _6906_ (.A(net426),
    .B(net245),
    .X(_3512_));
 sky130_fd_sc_hd__o211a_1 _6907_ (.A1(net3),
    .A2(net257),
    .B1(net165),
    .C1(_3512_),
    .X(_1195_));
 sky130_fd_sc_hd__nand2_1 _6908_ (.A(_1279_),
    .B(net259),
    .Y(_3513_));
 sky130_fd_sc_hd__o211a_1 _6909_ (.A1(net4),
    .A2(net259),
    .B1(net167),
    .C1(_3513_),
    .X(_1196_));
 sky130_fd_sc_hd__nand2_1 _6910_ (.A(_1278_),
    .B(net260),
    .Y(_3514_));
 sky130_fd_sc_hd__o211a_1 _6911_ (.A1(net5),
    .A2(net260),
    .B1(net167),
    .C1(_3514_),
    .X(_1197_));
 sky130_fd_sc_hd__or2_1 _6912_ (.A(net425),
    .B(net253),
    .X(_3515_));
 sky130_fd_sc_hd__o211a_1 _6913_ (.A1(net6),
    .A2(net264),
    .B1(net169),
    .C1(_3515_),
    .X(_1198_));
 sky130_fd_sc_hd__or2_1 _6914_ (.A(net408),
    .B(net248),
    .X(_3516_));
 sky130_fd_sc_hd__o211a_1 _6915_ (.A1(net7),
    .A2(net258),
    .B1(net166),
    .C1(_3516_),
    .X(_1199_));
 sky130_fd_sc_hd__or2_1 _6916_ (.A(net400),
    .B(net246),
    .X(_3517_));
 sky130_fd_sc_hd__o211a_1 _6917_ (.A1(net8),
    .A2(net255),
    .B1(net164),
    .C1(_3517_),
    .X(_1200_));
 sky130_fd_sc_hd__or2_1 _6918_ (.A(net399),
    .B(net244),
    .X(_3518_));
 sky130_fd_sc_hd__o211a_1 _6919_ (.A1(net9),
    .A2(net254),
    .B1(net165),
    .C1(_3518_),
    .X(_1201_));
 sky130_fd_sc_hd__or2_1 _6920_ (.A(net2020),
    .B(net253),
    .X(_3519_));
 sky130_fd_sc_hd__o211a_1 _6921_ (.A1(net10),
    .A2(net264),
    .B1(net169),
    .C1(_3519_),
    .X(_1202_));
 sky130_fd_sc_hd__or2_1 _6922_ (.A(net395),
    .B(net253),
    .X(_3520_));
 sky130_fd_sc_hd__o211a_1 _6923_ (.A1(net11),
    .A2(net264),
    .B1(net169),
    .C1(_3520_),
    .X(_1203_));
 sky130_fd_sc_hd__or2_1 _6924_ (.A(net378),
    .B(net248),
    .X(_3521_));
 sky130_fd_sc_hd__o211a_1 _6925_ (.A1(net12),
    .A2(net258),
    .B1(net166),
    .C1(_3521_),
    .X(_1204_));
 sky130_fd_sc_hd__or2_1 _6926_ (.A(net374),
    .B(net253),
    .X(_3522_));
 sky130_fd_sc_hd__o211a_1 _6927_ (.A1(net13),
    .A2(net264),
    .B1(net169),
    .C1(_3522_),
    .X(_1205_));
 sky130_fd_sc_hd__or2_1 _6928_ (.A(net368),
    .B(net248),
    .X(_3523_));
 sky130_fd_sc_hd__o211a_1 _6929_ (.A1(net14),
    .A2(net257),
    .B1(net164),
    .C1(_3523_),
    .X(_1206_));
 sky130_fd_sc_hd__or2_1 _6930_ (.A(net2221),
    .B(net250),
    .X(_3524_));
 sky130_fd_sc_hd__o211a_1 _6931_ (.A1(net15),
    .A2(net261),
    .B1(net170),
    .C1(_3524_),
    .X(_1207_));
 sky130_fd_sc_hd__or2_1 _6932_ (.A(net708),
    .B(net248),
    .X(_3525_));
 sky130_fd_sc_hd__o211a_1 _6933_ (.A1(net16),
    .A2(net258),
    .B1(net166),
    .C1(_3525_),
    .X(_1208_));
 sky130_fd_sc_hd__or2_1 _6934_ (.A(net2056),
    .B(net244),
    .X(_3526_));
 sky130_fd_sc_hd__o211a_1 _6935_ (.A1(net17),
    .A2(net254),
    .B1(net165),
    .C1(_3526_),
    .X(_1209_));
 sky130_fd_sc_hd__or2_1 _6936_ (.A(net587),
    .B(net253),
    .X(_3527_));
 sky130_fd_sc_hd__o211a_1 _6937_ (.A1(net18),
    .A2(net264),
    .B1(net169),
    .C1(_3527_),
    .X(_1210_));
 sky130_fd_sc_hd__or2_1 _6938_ (.A(net1924),
    .B(net244),
    .X(_3528_));
 sky130_fd_sc_hd__o211a_1 _6939_ (.A1(net19),
    .A2(net254),
    .B1(net165),
    .C1(_3528_),
    .X(_1211_));
 sky130_fd_sc_hd__or2_1 _6940_ (.A(net2106),
    .B(net253),
    .X(_3529_));
 sky130_fd_sc_hd__o211a_1 _6941_ (.A1(net20),
    .A2(net264),
    .B1(net169),
    .C1(_3529_),
    .X(_1212_));
 sky130_fd_sc_hd__or2_1 _6942_ (.A(net2018),
    .B(net247),
    .X(_3530_));
 sky130_fd_sc_hd__o211a_1 _6943_ (.A1(net22),
    .A2(net256),
    .B1(net164),
    .C1(_3530_),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_1 _6944_ (.A(_1277_),
    .B(net258),
    .Y(_3531_));
 sky130_fd_sc_hd__o211a_1 _6945_ (.A1(net23),
    .A2(net258),
    .B1(net166),
    .C1(_3531_),
    .X(_1214_));
 sky130_fd_sc_hd__mux2_1 _6946_ (.A0(net2082),
    .A1(net873),
    .S(net264),
    .X(_3532_));
 sky130_fd_sc_hd__nand2b_1 _6947_ (.A_N(_3532_),
    .B(net169),
    .Y(_1215_));
 sky130_fd_sc_hd__or2_1 _6948_ (.A(net839),
    .B(net252),
    .X(_3533_));
 sky130_fd_sc_hd__o211a_1 _6949_ (.A1(net2040),
    .A2(net263),
    .B1(net168),
    .C1(_3533_),
    .X(_1216_));
 sky130_fd_sc_hd__or2_1 _6950_ (.A(net628),
    .B(net252),
    .X(_3534_));
 sky130_fd_sc_hd__o211a_1 _6951_ (.A1(net2015),
    .A2(net263),
    .B1(net168),
    .C1(_3534_),
    .X(_1217_));
 sky130_fd_sc_hd__or2_1 _6952_ (.A(net606),
    .B(net251),
    .X(_3535_));
 sky130_fd_sc_hd__o211a_1 _6953_ (.A1(net2008),
    .A2(net262),
    .B1(net168),
    .C1(_3535_),
    .X(_1218_));
 sky130_fd_sc_hd__or2_1 _6954_ (.A(net551),
    .B(net250),
    .X(_3536_));
 sky130_fd_sc_hd__o211a_1 _6955_ (.A1(net1998),
    .A2(net260),
    .B1(net167),
    .C1(_3536_),
    .X(_1219_));
 sky130_fd_sc_hd__or2_1 _6956_ (.A(net875),
    .B(net249),
    .X(_3537_));
 sky130_fd_sc_hd__o211a_1 _6957_ (.A1(net949),
    .A2(net259),
    .B1(net167),
    .C1(_3537_),
    .X(_1220_));
 sky130_fd_sc_hd__or2_1 _6958_ (.A(net778),
    .B(net249),
    .X(_3538_));
 sky130_fd_sc_hd__o211a_1 _6959_ (.A1(net2017),
    .A2(net259),
    .B1(net167),
    .C1(_3538_),
    .X(_1221_));
 sky130_fd_sc_hd__or2_1 _6960_ (.A(net814),
    .B(net252),
    .X(_3539_));
 sky130_fd_sc_hd__o211a_1 _6961_ (.A1(net2016),
    .A2(net263),
    .B1(net168),
    .C1(_3539_),
    .X(_1222_));
 sky130_fd_sc_hd__or2_1 _6962_ (.A(net754),
    .B(net248),
    .X(_3540_));
 sky130_fd_sc_hd__o211a_1 _6963_ (.A1(net2043),
    .A2(net258),
    .B1(net166),
    .C1(_3540_),
    .X(_1223_));
 sky130_fd_sc_hd__or2_1 _6964_ (.A(net539),
    .B(net248),
    .X(_3541_));
 sky130_fd_sc_hd__o211a_1 _6965_ (.A1(net2065),
    .A2(net258),
    .B1(net166),
    .C1(_3541_),
    .X(_1224_));
 sky130_fd_sc_hd__or2_1 _6966_ (.A(net830),
    .B(net251),
    .X(_3542_));
 sky130_fd_sc_hd__o211a_1 _6967_ (.A1(net1741),
    .A2(net262),
    .B1(net168),
    .C1(_3542_),
    .X(_1225_));
 sky130_fd_sc_hd__or2_1 _6968_ (.A(net559),
    .B(net249),
    .X(_3543_));
 sky130_fd_sc_hd__o211a_1 _6969_ (.A1(net2027),
    .A2(net259),
    .B1(net167),
    .C1(_3543_),
    .X(_1226_));
 sky130_fd_sc_hd__or2_1 _6970_ (.A(net847),
    .B(net251),
    .X(_3544_));
 sky130_fd_sc_hd__o211a_1 _6971_ (.A1(net2009),
    .A2(net262),
    .B1(net168),
    .C1(_3544_),
    .X(_1227_));
 sky130_fd_sc_hd__or2_1 _6972_ (.A(net856),
    .B(net251),
    .X(_3545_));
 sky130_fd_sc_hd__o211a_1 _6973_ (.A1(net2083),
    .A2(net262),
    .B1(net168),
    .C1(_3545_),
    .X(_1228_));
 sky130_fd_sc_hd__or2_1 _6974_ (.A(net802),
    .B(net250),
    .X(_3546_));
 sky130_fd_sc_hd__o211a_1 _6975_ (.A1(net2062),
    .A2(net260),
    .B1(net167),
    .C1(_3546_),
    .X(_1229_));
 sky130_fd_sc_hd__or2_1 _6976_ (.A(net793),
    .B(net250),
    .X(_3547_));
 sky130_fd_sc_hd__o211a_1 _6977_ (.A1(net2034),
    .A2(net259),
    .B1(net167),
    .C1(_3547_),
    .X(_1230_));
 sky130_fd_sc_hd__or2_1 _6978_ (.A(net758),
    .B(net252),
    .X(_3548_));
 sky130_fd_sc_hd__o211a_1 _6979_ (.A1(net889),
    .A2(net263),
    .B1(net168),
    .C1(_3548_),
    .X(_1231_));
 sky130_fd_sc_hd__or2_1 _6980_ (.A(net718),
    .B(net248),
    .X(_3549_));
 sky130_fd_sc_hd__o211a_1 _6981_ (.A1(net2049),
    .A2(net258),
    .B1(net166),
    .C1(_3549_),
    .X(_1232_));
 sky130_fd_sc_hd__or2_1 _6982_ (.A(net810),
    .B(net246),
    .X(_3550_));
 sky130_fd_sc_hd__o211a_1 _6983_ (.A1(net2007),
    .A2(net255),
    .B1(net164),
    .C1(_3550_),
    .X(_1233_));
 sky130_fd_sc_hd__or2_1 _6984_ (.A(net656),
    .B(net246),
    .X(_3551_));
 sky130_fd_sc_hd__o211a_1 _6985_ (.A1(net2033),
    .A2(net255),
    .B1(net164),
    .C1(_3551_),
    .X(_1234_));
 sky130_fd_sc_hd__or2_1 _6986_ (.A(net863),
    .B(net244),
    .X(_3552_));
 sky130_fd_sc_hd__o211a_1 _6987_ (.A1(net2060),
    .A2(net254),
    .B1(net165),
    .C1(_3552_),
    .X(_1235_));
 sky130_fd_sc_hd__or2_1 _6988_ (.A(net861),
    .B(net246),
    .X(_3553_));
 sky130_fd_sc_hd__o211a_1 _6989_ (.A1(net2073),
    .A2(net255),
    .B1(net164),
    .C1(_3553_),
    .X(_1236_));
 sky130_fd_sc_hd__or2_1 _6990_ (.A(net2053),
    .B(net246),
    .X(_3554_));
 sky130_fd_sc_hd__o211a_1 _6991_ (.A1(net2047),
    .A2(net255),
    .B1(net164),
    .C1(_3554_),
    .X(_1237_));
 sky130_fd_sc_hd__or2_1 _6992_ (.A(net824),
    .B(net246),
    .X(_3555_));
 sky130_fd_sc_hd__o211a_1 _6993_ (.A1(net2036),
    .A2(net255),
    .B1(net164),
    .C1(_3555_),
    .X(_1238_));
 sky130_fd_sc_hd__or2_1 _6994_ (.A(net858),
    .B(net247),
    .X(_3556_));
 sky130_fd_sc_hd__o211a_1 _6995_ (.A1(net1955),
    .A2(net256),
    .B1(net164),
    .C1(_3556_),
    .X(_1239_));
 sky130_fd_sc_hd__or2_1 _6996_ (.A(net611),
    .B(net247),
    .X(_3557_));
 sky130_fd_sc_hd__o211a_1 _6997_ (.A1(net2066),
    .A2(net256),
    .B1(net164),
    .C1(_3557_),
    .X(_1240_));
 sky130_fd_sc_hd__or2_1 _6998_ (.A(net742),
    .B(net244),
    .X(_3558_));
 sky130_fd_sc_hd__o211a_1 _6999_ (.A1(net2025),
    .A2(net254),
    .B1(net165),
    .C1(_3558_),
    .X(_1241_));
 sky130_fd_sc_hd__or2_1 _7000_ (.A(net837),
    .B(net244),
    .X(_3559_));
 sky130_fd_sc_hd__o211a_1 _7001_ (.A1(net2051),
    .A2(net254),
    .B1(net165),
    .C1(_3559_),
    .X(_1242_));
 sky130_fd_sc_hd__or2_1 _7002_ (.A(net798),
    .B(net245),
    .X(_3560_));
 sky130_fd_sc_hd__o211a_1 _7003_ (.A1(net2061),
    .A2(net257),
    .B1(net165),
    .C1(_3560_),
    .X(_1243_));
 sky130_fd_sc_hd__or2_1 _7004_ (.A(net565),
    .B(net247),
    .X(_3561_));
 sky130_fd_sc_hd__o211a_1 _7005_ (.A1(net2041),
    .A2(net256),
    .B1(net164),
    .C1(_3561_),
    .X(_1244_));
 sky130_fd_sc_hd__and2_1 _7006_ (.A(net449),
    .B(net706),
    .X(_1275_));
 sky130_fd_sc_hd__and2_1 _7007_ (.A(net449),
    .B(net700),
    .X(_1276_));
 sky130_fd_sc_hd__o211a_1 _7008_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .A2(_2037_),
    .B1(_2035_),
    .C1(_2033_),
    .X(_3563_));
 sky130_fd_sc_hd__o211a_1 _7009_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .A2(_2037_),
    .B1(_2035_),
    .C1(_2033_),
    .X(_3564_));
 sky130_fd_sc_hd__o211a_1 _7010_ (.A1(net2247),
    .A2(_2037_),
    .B1(_2035_),
    .C1(_2033_),
    .X(_3565_));
 sky130_fd_sc_hd__o211a_1 _7011_ (.A1(net2029),
    .A2(_2037_),
    .B1(_2035_),
    .C1(_2033_),
    .X(_3566_));
 sky130_fd_sc_hd__inv_2 _7012_ (.A(net462),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _7013_ (.A(net461),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _7014_ (.A(net461),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _7015_ (.A(net461),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _7016_ (.A(net460),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _7017_ (.A(net460),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _7018_ (.A(net461),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _7019_ (.A(net461),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _7020_ (.A(net461),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _7021_ (.A(net461),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _7022_ (.A(net461),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _7023_ (.A(net461),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _7024_ (.A(net461),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _7025_ (.A(net462),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _7026_ (.A(net462),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _7027_ (.A(net462),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _7028_ (.A(net465),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _7029_ (.A(net458),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _7030_ (.A(net458),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _7031_ (.A(net457),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _7032_ (.A(net458),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _7033_ (.A(net458),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _7034_ (.A(net458),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _7035_ (.A(net458),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _7036_ (.A(net458),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _7037_ (.A(net457),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _7038_ (.A(net457),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _7039_ (.A(net459),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _7040_ (.A(net459),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _7041__2 (.A(clknet_leaf_36_clk),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _7042__3 (.A(clknet_leaf_35_clk),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _7043__4 (.A(clknet_leaf_32_clk),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _7044__5 (.A(clknet_leaf_25_clk),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _7045__6 (.A(clknet_leaf_23_clk),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _7046__7 (.A(clknet_leaf_52_clk),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _7047__8 (.A(clknet_leaf_42_clk),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _7048__9 (.A(clknet_leaf_44_clk),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _7049__10 (.A(clknet_leaf_29_clk),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _7050__11 (.A(clknet_leaf_47_clk),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _7051__12 (.A(clknet_leaf_70_clk),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _7052__13 (.A(clknet_leaf_23_clk),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _7053__14 (.A(clknet_leaf_51_clk),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _7054__15 (.A(clknet_leaf_22_clk),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _7055__16 (.A(clknet_leaf_18_clk),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _7056__17 (.A(clknet_leaf_40_clk),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _7057__18 (.A(clknet_leaf_19_clk),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _7058__19 (.A(clknet_leaf_27_clk),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _7059__20 (.A(clknet_leaf_47_clk),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _7060__21 (.A(clknet_leaf_72_clk),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _7061__22 (.A(clknet_leaf_55_clk),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _7062__23 (.A(clknet_leaf_38_clk),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _7063__24 (.A(clknet_leaf_58_clk),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _7064__25 (.A(clknet_leaf_26_clk),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _7065__26 (.A(clknet_leaf_64_clk),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _7066__27 (.A(clknet_leaf_58_clk),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _7067__28 (.A(clknet_leaf_51_clk),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _7068__29 (.A(clknet_leaf_78_clk),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _7069__30 (.A(clknet_leaf_71_clk),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _7070__31 (.A(clknet_leaf_56_clk),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _7071__32 (.A(clknet_leaf_56_clk),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _7072__33 (.A(clknet_leaf_33_clk),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _7073__34 (.A(clknet_leaf_36_clk),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _7074__35 (.A(clknet_leaf_35_clk),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _7075__36 (.A(clknet_leaf_32_clk),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _7076__37 (.A(clknet_leaf_25_clk),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _7077__38 (.A(clknet_leaf_23_clk),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _7078__39 (.A(clknet_leaf_51_clk),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _7079__40 (.A(clknet_leaf_42_clk),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _7080__41 (.A(clknet_leaf_45_clk),
    .Y(net513));
 sky130_fd_sc_hd__inv_2 _7081__42 (.A(clknet_leaf_30_clk),
    .Y(net514));
 sky130_fd_sc_hd__inv_2 _7082__43 (.A(clknet_leaf_47_clk),
    .Y(net515));
 sky130_fd_sc_hd__inv_2 _7083__44 (.A(clknet_leaf_70_clk),
    .Y(net516));
 sky130_fd_sc_hd__inv_2 _7084__45 (.A(clknet_leaf_23_clk),
    .Y(net517));
 sky130_fd_sc_hd__inv_2 _7085__46 (.A(clknet_leaf_52_clk),
    .Y(net518));
 sky130_fd_sc_hd__inv_2 _7086__47 (.A(clknet_leaf_21_clk),
    .Y(net519));
 sky130_fd_sc_hd__inv_2 _7087__48 (.A(clknet_leaf_14_clk),
    .Y(net520));
 sky130_fd_sc_hd__inv_2 _7088__49 (.A(clknet_leaf_40_clk),
    .Y(net521));
 sky130_fd_sc_hd__inv_2 _7089__50 (.A(clknet_leaf_20_clk),
    .Y(net522));
 sky130_fd_sc_hd__inv_2 _7090__51 (.A(clknet_leaf_26_clk),
    .Y(net523));
 sky130_fd_sc_hd__inv_2 _7091__52 (.A(clknet_leaf_51_clk),
    .Y(net524));
 sky130_fd_sc_hd__inv_2 _7092__53 (.A(clknet_leaf_72_clk),
    .Y(net525));
 sky130_fd_sc_hd__inv_2 _7093__54 (.A(clknet_leaf_55_clk),
    .Y(net526));
 sky130_fd_sc_hd__inv_2 _7094__55 (.A(clknet_leaf_38_clk),
    .Y(net527));
 sky130_fd_sc_hd__inv_2 _7095__56 (.A(clknet_leaf_58_clk),
    .Y(net528));
 sky130_fd_sc_hd__inv_2 _7096__57 (.A(clknet_leaf_29_clk),
    .Y(net529));
 sky130_fd_sc_hd__inv_2 _7097__58 (.A(clknet_leaf_64_clk),
    .Y(net530));
 sky130_fd_sc_hd__inv_2 _7098__59 (.A(clknet_leaf_59_clk),
    .Y(net531));
 sky130_fd_sc_hd__inv_2 _7099__60 (.A(clknet_leaf_52_clk),
    .Y(net532));
 sky130_fd_sc_hd__inv_2 _7100__61 (.A(clknet_leaf_70_clk),
    .Y(net533));
 sky130_fd_sc_hd__inv_2 _7101__62 (.A(clknet_leaf_71_clk),
    .Y(net534));
 sky130_fd_sc_hd__inv_2 _7102__63 (.A(clknet_leaf_50_clk),
    .Y(net535));
 sky130_fd_sc_hd__inv_2 _7103__64 (.A(clknet_leaf_55_clk),
    .Y(net536));
 sky130_fd_sc_hd__inv_2 _7104_ (.A(net465),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _7105_ (.A(net462),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _7106_ (.A(net461),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _7107_ (.A(net461),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _7108_ (.A(net462),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _7109_ (.A(net460),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _7110_ (.A(net460),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _7111_ (.A(net463),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _7112_ (.A(net63),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _7113_ (.A(net461),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _7114_ (.A(net463),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _7115_ (.A(net465),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _7116_ (.A(net463),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _7117_ (.A(net462),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _7118_ (.A(net460),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _7119_ (.A(net462),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _7120_ (.A(net463),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _7121_ (.A(net465),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _7122_ (.A(net458),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _7123_ (.A(net458),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _7124_ (.A(net457),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _7125_ (.A(net457),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _7126_ (.A(net458),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _7127_ (.A(net458),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _7128_ (.A(net459),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _7129_ (.A(net457),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _7130_ (.A(net457),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _7131_ (.A(net457),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _7132_ (.A(net459),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _7133_ (.A(net459),
    .Y(_0192_));
 sky130_fd_sc_hd__dfxtp_1 _7134_ (.CLK(clknet_leaf_78_clk),
    .D(_0193_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7135_ (.CLK(clknet_leaf_79_clk),
    .D(_0194_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7136_ (.CLK(clknet_leaf_78_clk),
    .D(_0195_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7137_ (.CLK(clknet_leaf_78_clk),
    .D(_0196_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ));
 sky130_fd_sc_hd__dfxtp_2 _7138_ (.CLK(clknet_leaf_45_clk),
    .D(net589),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7139_ (.CLK(clknet_leaf_68_clk),
    .D(_0198_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7140_ (.CLK(clknet_leaf_76_clk),
    .D(_0199_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ));
 sky130_fd_sc_hd__dfxtp_2 _7141_ (.CLK(clknet_leaf_45_clk),
    .D(net580),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7142_ (.CLK(clknet_leaf_72_clk),
    .D(net1191),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7143_ (.CLK(clknet_leaf_69_clk),
    .D(_0202_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7144_ (.CLK(clknet_leaf_71_clk),
    .D(net922),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7145_ (.CLK(clknet_leaf_65_clk),
    .D(net1716),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7146_ (.CLK(clknet_leaf_44_clk),
    .D(net2022),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7147_ (.CLK(clknet_leaf_44_clk),
    .D(_0206_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7148_ (.CLK(clknet_leaf_46_clk),
    .D(_0207_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7149_ (.CLK(clknet_leaf_17_clk),
    .D(_0208_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7150_ (.CLK(clknet_leaf_17_clk),
    .D(_0209_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7151_ (.CLK(clknet_leaf_3_clk),
    .D(_0210_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7152_ (.CLK(clknet_leaf_3_clk),
    .D(_0211_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7153_ (.CLK(clknet_leaf_15_clk),
    .D(_0212_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ));
 sky130_fd_sc_hd__dfxtp_2 _7154_ (.CLK(clknet_leaf_4_clk),
    .D(net2031),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7155_ (.CLK(clknet_leaf_2_clk),
    .D(_0214_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7156_ (.CLK(clknet_leaf_15_clk),
    .D(_0215_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7157_ (.CLK(clknet_leaf_3_clk),
    .D(net2039),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7158_ (.CLK(clknet_leaf_15_clk),
    .D(_0217_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7159_ (.CLK(clknet_leaf_15_clk),
    .D(_0218_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7160_ (.CLK(clknet_leaf_15_clk),
    .D(net709),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7161_ (.CLK(clknet_leaf_17_clk),
    .D(_0220_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7162_ (.CLK(clknet_leaf_17_clk),
    .D(_0221_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7163_ (.CLK(clknet_leaf_18_clk),
    .D(_0222_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7164_ (.CLK(clknet_leaf_17_clk),
    .D(_0223_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7165_ (.CLK(clknet_leaf_3_clk),
    .D(_0224_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7166_ (.CLK(clknet_leaf_1_clk),
    .D(_0225_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7167_ (.CLK(clknet_leaf_1_clk),
    .D(_0226_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7168_ (.CLK(clknet_leaf_1_clk),
    .D(_0227_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7169_ (.CLK(clknet_leaf_13_clk),
    .D(_0228_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7170_ (.CLK(clknet_leaf_33_clk),
    .D(net2097),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7171_ (.CLK(clknet_leaf_36_clk),
    .D(net1837),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7172_ (.CLK(clknet_leaf_36_clk),
    .D(net1883),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7173_ (.CLK(clknet_leaf_32_clk),
    .D(net1903),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7174_ (.CLK(clknet_leaf_24_clk),
    .D(net1833),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7175_ (.CLK(clknet_leaf_24_clk),
    .D(net1806),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7176_ (.CLK(clknet_leaf_53_clk),
    .D(net1646),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7177_ (.CLK(clknet_leaf_42_clk),
    .D(net1839),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7178_ (.CLK(clknet_leaf_41_clk),
    .D(net1877),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7179_ (.CLK(clknet_leaf_30_clk),
    .D(net1747),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7180_ (.CLK(clknet_leaf_51_clk),
    .D(net2002),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7181_ (.CLK(clknet_leaf_69_clk),
    .D(net1764),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7182_ (.CLK(clknet_leaf_23_clk),
    .D(net1989),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7183_ (.CLK(clknet_leaf_53_clk),
    .D(net1718),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7184_ (.CLK(clknet_leaf_23_clk),
    .D(net1943),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7185_ (.CLK(clknet_leaf_22_clk),
    .D(net1669),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7186_ (.CLK(clknet_leaf_39_clk),
    .D(net1760),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7187_ (.CLK(clknet_leaf_20_clk),
    .D(net1788),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7188_ (.CLK(clknet_leaf_26_clk),
    .D(net1871),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(clknet_leaf_51_clk),
    .D(net1935),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(clknet_leaf_72_clk),
    .D(net1766),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7191_ (.CLK(clknet_leaf_55_clk),
    .D(net1817),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(clknet_leaf_38_clk),
    .D(net1753),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7193_ (.CLK(clknet_leaf_60_clk),
    .D(net1865),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(clknet_leaf_30_clk),
    .D(net1786),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(clknet_leaf_63_clk),
    .D(net1745),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(clknet_leaf_60_clk),
    .D(net1671),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7197_ (.CLK(clknet_leaf_53_clk),
    .D(net1614),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7198_ (.CLK(clknet_leaf_70_clk),
    .D(net1891),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7199_ (.CLK(clknet_leaf_64_clk),
    .D(net1808),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7200_ (.CLK(clknet_leaf_49_clk),
    .D(net1652),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7201_ (.CLK(clknet_leaf_59_clk),
    .D(net1778),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7202_ (.CLK(clknet_leaf_33_clk),
    .D(net1770),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7203_ (.CLK(clknet_leaf_36_clk),
    .D(net2094),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7204_ (.CLK(clknet_leaf_42_clk),
    .D(net1907),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7205_ (.CLK(clknet_leaf_32_clk),
    .D(net1815),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7206_ (.CLK(clknet_leaf_24_clk),
    .D(net1869),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7207_ (.CLK(clknet_leaf_24_clk),
    .D(net1804),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7208_ (.CLK(clknet_leaf_52_clk),
    .D(net1798),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7209_ (.CLK(clknet_leaf_42_clk),
    .D(net1921),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7210_ (.CLK(clknet_leaf_45_clk),
    .D(net1847),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7211_ (.CLK(clknet_leaf_30_clk),
    .D(net1738),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7212_ (.CLK(clknet_leaf_51_clk),
    .D(net1991),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7213_ (.CLK(clknet_leaf_69_clk),
    .D(net1813),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7214_ (.CLK(clknet_leaf_24_clk),
    .D(net1849),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7215_ (.CLK(clknet_leaf_54_clk),
    .D(net1897),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7216_ (.CLK(clknet_leaf_22_clk),
    .D(net1913),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7217_ (.CLK(clknet_leaf_18_clk),
    .D(net1843),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7218_ (.CLK(clknet_leaf_40_clk),
    .D(net1881),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7219_ (.CLK(clknet_leaf_19_clk),
    .D(net1855),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7220_ (.CLK(clknet_leaf_25_clk),
    .D(net1827),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7221_ (.CLK(clknet_leaf_47_clk),
    .D(net1905),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7222_ (.CLK(clknet_leaf_72_clk),
    .D(net1774),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7223_ (.CLK(clknet_leaf_55_clk),
    .D(net1821),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7224_ (.CLK(clknet_leaf_38_clk),
    .D(net1768),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7225_ (.CLK(clknet_leaf_63_clk),
    .D(net1755),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7226_ (.CLK(clknet_leaf_26_clk),
    .D(net1873),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7227_ (.CLK(clknet_leaf_64_clk),
    .D(net1950),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7228_ (.CLK(clknet_leaf_60_clk),
    .D(net1819),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7229_ (.CLK(clknet_leaf_52_clk),
    .D(net1845),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7230_ (.CLK(clknet_leaf_69_clk),
    .D(net1810),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7231_ (.CLK(clknet_leaf_65_clk),
    .D(net1728),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7232_ (.CLK(clknet_leaf_49_clk),
    .D(net1706),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7233_ (.CLK(clknet_leaf_59_clk),
    .D(net1612),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ));
 sky130_fd_sc_hd__dfstp_1 _7234_ (.CLK(clknet_leaf_20_clk),
    .D(_0293_),
    .SET_B(net453),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7235_ (.CLK(clknet_leaf_14_clk),
    .D(_0294_),
    .RESET_B(_0070_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7236_ (.CLK(clknet_leaf_14_clk),
    .D(_0295_),
    .RESET_B(_0071_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7237_ (.CLK(clknet_leaf_14_clk),
    .D(_0296_),
    .RESET_B(_0072_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7238_ (.CLK(clknet_leaf_14_clk),
    .D(_0297_),
    .RESET_B(_0073_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7239_ (.CLK(clknet_leaf_5_clk),
    .D(_0298_),
    .RESET_B(_0074_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7240_ (.CLK(clknet_leaf_5_clk),
    .D(_0299_),
    .RESET_B(_0075_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7241_ (.CLK(clknet_leaf_13_clk),
    .D(_0300_),
    .RESET_B(_0076_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7242_ (.CLK(clknet_leaf_13_clk),
    .D(_0301_),
    .RESET_B(_0077_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7243_ (.CLK(clknet_leaf_13_clk),
    .D(_0302_),
    .RESET_B(_0078_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7244_ (.CLK(clknet_leaf_13_clk),
    .D(_0303_),
    .RESET_B(_0079_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7245_ (.CLK(clknet_leaf_13_clk),
    .D(_0304_),
    .RESET_B(_0080_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7246_ (.CLK(clknet_leaf_12_clk),
    .D(_0305_),
    .RESET_B(_0081_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7247_ (.CLK(clknet_leaf_13_clk),
    .D(_0306_),
    .RESET_B(_0082_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7248_ (.CLK(clknet_leaf_17_clk),
    .D(net2063),
    .RESET_B(_0083_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7249_ (.CLK(clknet_leaf_18_clk),
    .D(net2035),
    .RESET_B(_0084_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7250_ (.CLK(clknet_leaf_18_clk),
    .D(_0309_),
    .RESET_B(_0085_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7251_ (.CLK(clknet_leaf_47_clk),
    .D(_0310_),
    .RESET_B(_0086_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7252_ (.CLK(clknet_leaf_67_clk),
    .D(_0311_),
    .RESET_B(_0087_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7253_ (.CLK(clknet_leaf_67_clk),
    .D(_0312_),
    .RESET_B(_0088_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7254_ (.CLK(clknet_leaf_67_clk),
    .D(_0313_),
    .RESET_B(_0089_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7255_ (.CLK(clknet_leaf_66_clk),
    .D(net2074),
    .RESET_B(_0090_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7256_ (.CLK(clknet_leaf_66_clk),
    .D(net2048),
    .RESET_B(_0091_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7257_ (.CLK(clknet_leaf_66_clk),
    .D(_0316_),
    .RESET_B(_0092_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7258_ (.CLK(clknet_leaf_62_clk),
    .D(_0317_),
    .RESET_B(_0093_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7259_ (.CLK(clknet_leaf_62_clk),
    .D(_0318_),
    .RESET_B(_0094_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7260_ (.CLK(clknet_leaf_80_clk),
    .D(_0319_),
    .RESET_B(_0095_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7261_ (.CLK(clknet_leaf_79_clk),
    .D(_0320_),
    .RESET_B(_0096_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7262_ (.CLK(clknet_leaf_79_clk),
    .D(_0321_),
    .RESET_B(_0097_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7263_ (.CLK(clknet_leaf_62_clk),
    .D(_0322_),
    .RESET_B(_0098_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7264_ (.CLK(clknet_leaf_34_clk),
    .D(net1156),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7265_ (.CLK(clknet_leaf_34_clk),
    .D(net896),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7266_ (.CLK(clknet_leaf_35_clk),
    .D(net1132),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7267_ (.CLK(clknet_leaf_34_clk),
    .D(net1536),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7268_ (.CLK(clknet_leaf_25_clk),
    .D(net1118),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7269_ (.CLK(clknet_leaf_23_clk),
    .D(net1488),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7270_ (.CLK(clknet_leaf_51_clk),
    .D(net1654),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7271_ (.CLK(clknet_leaf_44_clk),
    .D(net1184),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7272_ (.CLK(clknet_leaf_44_clk),
    .D(net1319),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7273_ (.CLK(clknet_leaf_29_clk),
    .D(net1350),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7274_ (.CLK(clknet_leaf_47_clk),
    .D(net1494),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7275_ (.CLK(clknet_leaf_70_clk),
    .D(net1606),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7276_ (.CLK(clknet_leaf_23_clk),
    .D(net1484),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7277_ (.CLK(clknet_leaf_50_clk),
    .D(net1301),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7278_ (.CLK(clknet_leaf_21_clk),
    .D(net1182),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7279_ (.CLK(clknet_leaf_21_clk),
    .D(net1364),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7280_ (.CLK(clknet_leaf_40_clk),
    .D(net1556),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7281_ (.CLK(clknet_leaf_20_clk),
    .D(net1168),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7282_ (.CLK(clknet_leaf_27_clk),
    .D(net1474),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7283_ (.CLK(clknet_leaf_50_clk),
    .D(net1050),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7284_ (.CLK(clknet_leaf_48_clk),
    .D(net1436),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7285_ (.CLK(clknet_leaf_56_clk),
    .D(net1313),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7286_ (.CLK(clknet_leaf_40_clk),
    .D(net1195),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7287_ (.CLK(clknet_leaf_64_clk),
    .D(net1558),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7288_ (.CLK(clknet_leaf_29_clk),
    .D(net1508),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7289_ (.CLK(clknet_leaf_64_clk),
    .D(net1584),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7290_ (.CLK(clknet_leaf_58_clk),
    .D(net1354),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7291_ (.CLK(clknet_leaf_51_clk),
    .D(net1544),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7292_ (.CLK(clknet_leaf_70_clk),
    .D(net1580),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7293_ (.CLK(clknet_leaf_71_clk),
    .D(net1261),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7294_ (.CLK(clknet_leaf_50_clk),
    .D(net1138),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7295_ (.CLK(clknet_leaf_56_clk),
    .D(net1336),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7296_ (.CLK(clknet_leaf_32_clk),
    .D(net1927),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7297_ (.CLK(clknet_leaf_33_clk),
    .D(net1965),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7298_ (.CLK(clknet_leaf_35_clk),
    .D(net1841),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7299_ (.CLK(clknet_leaf_32_clk),
    .D(net2102),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7300_ (.CLK(clknet_leaf_25_clk),
    .D(net1895),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7301_ (.CLK(clknet_leaf_25_clk),
    .D(net1987),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7302_ (.CLK(clknet_leaf_52_clk),
    .D(net1917),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7303_ (.CLK(clknet_leaf_42_clk),
    .D(net1995),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7304_ (.CLK(clknet_leaf_42_clk),
    .D(net1954),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7305_ (.CLK(clknet_leaf_31_clk),
    .D(net1732),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7306_ (.CLK(clknet_leaf_41_clk),
    .D(net1909),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7307_ (.CLK(clknet_leaf_72_clk),
    .D(net1851),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7308_ (.CLK(clknet_leaf_25_clk),
    .D(net1968),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7309_ (.CLK(clknet_leaf_54_clk),
    .D(net1975),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7310_ (.CLK(clknet_leaf_20_clk),
    .D(net1933),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7311_ (.CLK(clknet_leaf_19_clk),
    .D(net1823),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7312_ (.CLK(clknet_leaf_39_clk),
    .D(net1784),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7313_ (.CLK(clknet_leaf_35_clk),
    .D(net1835),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7314_ (.CLK(clknet_leaf_26_clk),
    .D(net1981),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7315_ (.CLK(clknet_leaf_50_clk),
    .D(net1919),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7316_ (.CLK(clknet_leaf_48_clk),
    .D(net2000),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7317_ (.CLK(clknet_leaf_54_clk),
    .D(net1831),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7318_ (.CLK(clknet_leaf_38_clk),
    .D(net1941),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7319_ (.CLK(clknet_leaf_58_clk),
    .D(net1970),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7320_ (.CLK(clknet_leaf_30_clk),
    .D(net1952),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7321_ (.CLK(clknet_leaf_57_clk),
    .D(net1875),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7322_ (.CLK(clknet_leaf_59_clk),
    .D(net1929),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7323_ (.CLK(clknet_leaf_52_clk),
    .D(net1939),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7324_ (.CLK(clknet_leaf_71_clk),
    .D(net1740),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7325_ (.CLK(clknet_leaf_64_clk),
    .D(net1979),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7326_ (.CLK(clknet_leaf_56_clk),
    .D(net1993),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7327_ (.CLK(clknet_leaf_59_clk),
    .D(net1861),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7328_ (.CLK(clknet_leaf_33_clk),
    .D(net878),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7329_ (.CLK(clknet_leaf_34_clk),
    .D(net882),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7330_ (.CLK(clknet_leaf_35_clk),
    .D(net1052),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7331_ (.CLK(clknet_leaf_34_clk),
    .D(net1134),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7332_ (.CLK(clknet_leaf_27_clk),
    .D(net1681),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7333_ (.CLK(clknet_leaf_27_clk),
    .D(net1241),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7334_ (.CLK(clknet_leaf_52_clk),
    .D(net1468),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7335_ (.CLK(clknet_leaf_42_clk),
    .D(net1644),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7336_ (.CLK(clknet_leaf_44_clk),
    .D(net1271),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7337_ (.CLK(clknet_leaf_30_clk),
    .D(net1164),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7338_ (.CLK(clknet_leaf_45_clk),
    .D(net1223),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7339_ (.CLK(clknet_leaf_71_clk),
    .D(net1384),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7340_ (.CLK(clknet_leaf_25_clk),
    .D(net1305),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7341_ (.CLK(clknet_leaf_50_clk),
    .D(net1126),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7342_ (.CLK(clknet_leaf_20_clk),
    .D(net1219),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7343_ (.CLK(clknet_leaf_19_clk),
    .D(net1088),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7344_ (.CLK(clknet_leaf_40_clk),
    .D(net1665),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7345_ (.CLK(clknet_leaf_35_clk),
    .D(net1506),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7346_ (.CLK(clknet_leaf_26_clk),
    .D(net1259),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7347_ (.CLK(clknet_leaf_50_clk),
    .D(net1114),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7348_ (.CLK(clknet_leaf_48_clk),
    .D(net1675),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7349_ (.CLK(clknet_leaf_56_clk),
    .D(net1685),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7350_ (.CLK(clknet_leaf_40_clk),
    .D(net1596),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7351_ (.CLK(clknet_leaf_64_clk),
    .D(net1630),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7352_ (.CLK(clknet_leaf_29_clk),
    .D(net1388),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7353_ (.CLK(clknet_leaf_64_clk),
    .D(net1859),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7354_ (.CLK(clknet_leaf_58_clk),
    .D(net1166),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7355_ (.CLK(clknet_leaf_51_clk),
    .D(net1372),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7356_ (.CLK(clknet_leaf_70_clk),
    .D(net1578),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7357_ (.CLK(clknet_leaf_71_clk),
    .D(net1500),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7358_ (.CLK(clknet_leaf_50_clk),
    .D(net1042),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7359_ (.CLK(clknet_leaf_57_clk),
    .D(net1040),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7360_ (.CLK(clknet_leaf_36_clk),
    .D(net1985),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7361_ (.CLK(clknet_leaf_36_clk),
    .D(net1977),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7362_ (.CLK(clknet_leaf_36_clk),
    .D(net2112),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7363_ (.CLK(clknet_leaf_31_clk),
    .D(net1945),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7364_ (.CLK(clknet_leaf_25_clk),
    .D(net1983),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7365_ (.CLK(clknet_leaf_24_clk),
    .D(net1776),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7366_ (.CLK(clknet_leaf_53_clk),
    .D(net1693),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7367_ (.CLK(clknet_leaf_40_clk),
    .D(net1889),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7368_ (.CLK(clknet_leaf_45_clk),
    .D(net1972),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7369_ (.CLK(clknet_leaf_31_clk),
    .D(net1667),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7370_ (.CLK(clknet_leaf_40_clk),
    .D(net1937),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7371_ (.CLK(clknet_leaf_71_clk),
    .D(net1963),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7372_ (.CLK(clknet_leaf_24_clk),
    .D(net1863),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7373_ (.CLK(clknet_leaf_54_clk),
    .D(net1899),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7374_ (.CLK(clknet_leaf_21_clk),
    .D(net1762),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7375_ (.CLK(clknet_leaf_21_clk),
    .D(net1893),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7376_ (.CLK(clknet_leaf_39_clk),
    .D(net1879),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7377_ (.CLK(clknet_leaf_28_clk),
    .D(net1885),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7378_ (.CLK(clknet_leaf_30_clk),
    .D(net1825),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7379_ (.CLK(clknet_leaf_50_clk),
    .D(net1911),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7380_ (.CLK(clknet_leaf_49_clk),
    .D(net1790),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7381_ (.CLK(clknet_leaf_54_clk),
    .D(net1997),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7382_ (.CLK(clknet_leaf_37_clk),
    .D(net1853),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7383_ (.CLK(clknet_leaf_58_clk),
    .D(net1923),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7384_ (.CLK(clknet_leaf_30_clk),
    .D(net1792),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7385_ (.CLK(clknet_leaf_64_clk),
    .D(net1931),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7386_ (.CLK(clknet_leaf_59_clk),
    .D(net1857),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7387_ (.CLK(clknet_leaf_39_clk),
    .D(net1800),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7388_ (.CLK(clknet_leaf_71_clk),
    .D(net1772),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7389_ (.CLK(clknet_leaf_64_clk),
    .D(net1901),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7390_ (.CLK(clknet_leaf_56_clk),
    .D(net1961),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7391_ (.CLK(clknet_leaf_55_clk),
    .D(net1958),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7392_ (.CLK(clknet_leaf_33_clk),
    .D(net971),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7393_ (.CLK(clknet_leaf_33_clk),
    .D(net1720),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7394_ (.CLK(clknet_leaf_42_clk),
    .D(net1683),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7395_ (.CLK(clknet_leaf_32_clk),
    .D(net1058),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7396_ (.CLK(clknet_leaf_24_clk),
    .D(net1307),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7397_ (.CLK(clknet_leaf_24_clk),
    .D(net1150),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7398_ (.CLK(clknet_leaf_53_clk),
    .D(net984),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7399_ (.CLK(clknet_leaf_40_clk),
    .D(net1576),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7400_ (.CLK(clknet_leaf_45_clk),
    .D(net1460),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7401_ (.CLK(clknet_leaf_30_clk),
    .D(net1029),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7402_ (.CLK(clknet_leaf_51_clk),
    .D(net1462),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7403_ (.CLK(clknet_leaf_69_clk),
    .D(net1038),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7404_ (.CLK(clknet_leaf_23_clk),
    .D(net1472),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7405_ (.CLK(clknet_leaf_53_clk),
    .D(net1398),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7406_ (.CLK(clknet_leaf_22_clk),
    .D(net1098),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7407_ (.CLK(clknet_leaf_18_clk),
    .D(net1015),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7408_ (.CLK(clknet_leaf_38_clk),
    .D(net1297),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7409_ (.CLK(clknet_leaf_19_clk),
    .D(net1162),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7410_ (.CLK(clknet_leaf_25_clk),
    .D(net1122),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7411_ (.CLK(clknet_leaf_47_clk),
    .D(net1332),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7412_ (.CLK(clknet_leaf_72_clk),
    .D(net1072),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7413_ (.CLK(clknet_leaf_55_clk),
    .D(net1299),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7414_ (.CLK(clknet_leaf_38_clk),
    .D(net1396),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7415_ (.CLK(clknet_leaf_60_clk),
    .D(net1217),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7416_ (.CLK(clknet_leaf_26_clk),
    .D(net1146),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7417_ (.CLK(clknet_leaf_64_clk),
    .D(net1406),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7418_ (.CLK(clknet_leaf_60_clk),
    .D(net1730),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7419_ (.CLK(clknet_leaf_52_clk),
    .D(net1356),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7420_ (.CLK(clknet_leaf_70_clk),
    .D(net1247),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7421_ (.CLK(clknet_leaf_65_clk),
    .D(net962),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7422_ (.CLK(clknet_leaf_49_clk),
    .D(net986),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7423_ (.CLK(clknet_leaf_59_clk),
    .D(net1289),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7424_ (.CLK(net473),
    .D(_0032_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7425_ (.CLK(net474),
    .D(_0043_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7426_ (.CLK(net475),
    .D(_0054_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7427_ (.CLK(net476),
    .D(_0057_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7428_ (.CLK(net477),
    .D(_0058_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7429_ (.CLK(net478),
    .D(_0059_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7430_ (.CLK(net479),
    .D(_0060_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7431_ (.CLK(net480),
    .D(_0061_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7432_ (.CLK(net481),
    .D(_0062_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7433_ (.CLK(net482),
    .D(_0063_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7434_ (.CLK(net483),
    .D(_0033_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7435_ (.CLK(net484),
    .D(_0034_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7436_ (.CLK(net485),
    .D(_0035_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7437_ (.CLK(net486),
    .D(_0036_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7438_ (.CLK(net487),
    .D(_0037_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7439_ (.CLK(net488),
    .D(_0038_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7440_ (.CLK(net489),
    .D(_0039_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7441_ (.CLK(net490),
    .D(_0040_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7442_ (.CLK(net491),
    .D(_0041_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7443_ (.CLK(net492),
    .D(_0042_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7444_ (.CLK(net493),
    .D(_0044_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7445_ (.CLK(net494),
    .D(_0045_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7446_ (.CLK(net495),
    .D(_0046_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7447_ (.CLK(net496),
    .D(_0047_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7448_ (.CLK(net497),
    .D(_0048_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7449_ (.CLK(net498),
    .D(_0049_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7450_ (.CLK(net499),
    .D(_0050_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7451_ (.CLK(net500),
    .D(_0051_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7452_ (.CLK(net501),
    .D(_0052_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7453_ (.CLK(net502),
    .D(_0053_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7454_ (.CLK(net503),
    .D(_0055_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7455_ (.CLK(net504),
    .D(_0056_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7456_ (.CLK(clknet_leaf_1_clk),
    .D(_0483_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7457_ (.CLK(clknet_leaf_24_clk),
    .D(_0484_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7458_ (.CLK(clknet_leaf_9_clk),
    .D(_0485_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7459_ (.CLK(clknet_leaf_77_clk),
    .D(_0486_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7460_ (.CLK(clknet_leaf_37_clk),
    .D(_0487_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7461_ (.CLK(clknet_leaf_37_clk),
    .D(_0488_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7462_ (.CLK(clknet_leaf_35_clk),
    .D(_0489_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7463_ (.CLK(clknet_leaf_23_clk),
    .D(_0490_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7464_ (.CLK(clknet_leaf_10_clk),
    .D(_0491_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7465_ (.CLK(clknet_leaf_11_clk),
    .D(_0492_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7466_ (.CLK(clknet_leaf_41_clk),
    .D(_0493_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7467_ (.CLK(clknet_leaf_15_clk),
    .D(_0494_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7468_ (.CLK(clknet_leaf_3_clk),
    .D(_0495_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7469_ (.CLK(clknet_leaf_10_clk),
    .D(_0496_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7470_ (.CLK(clknet_leaf_77_clk),
    .D(_0497_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7471_ (.CLK(clknet_leaf_78_clk),
    .D(_0498_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7472_ (.CLK(clknet_leaf_11_clk),
    .D(_0499_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7473_ (.CLK(clknet_leaf_47_clk),
    .D(_0500_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7474_ (.CLK(clknet_leaf_11_clk),
    .D(_0501_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7475_ (.CLK(clknet_leaf_13_clk),
    .D(_0502_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7476_ (.CLK(clknet_leaf_45_clk),
    .D(_0503_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7477_ (.CLK(clknet_leaf_19_clk),
    .D(_0504_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7478_ (.CLK(clknet_leaf_27_clk),
    .D(_0505_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7479_ (.CLK(clknet_leaf_48_clk),
    .D(_0506_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7480_ (.CLK(clknet_leaf_64_clk),
    .D(_0507_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7481_ (.CLK(clknet_leaf_61_clk),
    .D(_0508_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7482_ (.CLK(clknet_leaf_67_clk),
    .D(_0509_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7483_ (.CLK(clknet_leaf_66_clk),
    .D(_0510_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7484_ (.CLK(clknet_leaf_48_clk),
    .D(_0511_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7485_ (.CLK(clknet_leaf_62_clk),
    .D(net538),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7486_ (.CLK(clknet_leaf_60_clk),
    .D(_0513_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7487_ (.CLK(clknet_leaf_54_clk),
    .D(_0514_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7488_ (.CLK(clknet_leaf_68_clk),
    .D(_0515_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7489_ (.CLK(clknet_leaf_78_clk),
    .D(_0516_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7490_ (.CLK(clknet_leaf_76_clk),
    .D(_0517_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7491_ (.CLK(clknet_leaf_60_clk),
    .D(_0518_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7492_ (.CLK(clknet_leaf_37_clk),
    .D(net1542),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7493_ (.CLK(clknet_leaf_36_clk),
    .D(net809),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7494_ (.CLK(clknet_leaf_28_clk),
    .D(net785),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7495_ (.CLK(clknet_leaf_10_clk),
    .D(net591),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7496_ (.CLK(clknet_leaf_10_clk),
    .D(net705),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7497_ (.CLK(clknet_leaf_11_clk),
    .D(net661),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7498_ (.CLK(clknet_leaf_43_clk),
    .D(net641),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7499_ (.CLK(clknet_leaf_15_clk),
    .D(net633),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7500_ (.CLK(clknet_leaf_5_clk),
    .D(net745),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7501_ (.CLK(clknet_leaf_10_clk),
    .D(net781),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7502_ (.CLK(clknet_leaf_77_clk),
    .D(net593),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7503_ (.CLK(clknet_leaf_78_clk),
    .D(net721),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7504_ (.CLK(clknet_leaf_12_clk),
    .D(net739),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7505_ (.CLK(clknet_leaf_47_clk),
    .D(net601),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7506_ (.CLK(clknet_leaf_11_clk),
    .D(net725),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7507_ (.CLK(clknet_leaf_13_clk),
    .D(net763),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7508_ (.CLK(clknet_leaf_46_clk),
    .D(net554),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7509_ (.CLK(clknet_leaf_19_clk),
    .D(net649),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7510_ (.CLK(clknet_leaf_27_clk),
    .D(net681),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7511_ (.CLK(clknet_leaf_48_clk),
    .D(net691),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7512_ (.CLK(clknet_leaf_65_clk),
    .D(net620),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7513_ (.CLK(clknet_leaf_61_clk),
    .D(net603),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7514_ (.CLK(clknet_leaf_69_clk),
    .D(net790),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7515_ (.CLK(clknet_leaf_65_clk),
    .D(net663),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7516_ (.CLK(clknet_leaf_65_clk),
    .D(net637),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7517_ (.CLK(clknet_leaf_62_clk),
    .D(net655),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7518_ (.CLK(clknet_leaf_60_clk),
    .D(net570),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7519_ (.CLK(clknet_leaf_55_clk),
    .D(net958),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7520_ (.CLK(clknet_leaf_68_clk),
    .D(net639),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7521_ (.CLK(clknet_leaf_78_clk),
    .D(net599),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7522_ (.CLK(clknet_leaf_79_clk),
    .D(net749),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7523_ (.CLK(clknet_leaf_60_clk),
    .D(net715),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7524_ (.CLK(clknet_leaf_28_clk),
    .D(net624),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7525_ (.CLK(clknet_leaf_10_clk),
    .D(net574),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7526_ (.CLK(clknet_leaf_10_clk),
    .D(net761),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7527_ (.CLK(clknet_leaf_11_clk),
    .D(net687),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7528_ (.CLK(clknet_leaf_43_clk),
    .D(net665),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7529_ (.CLK(clknet_leaf_15_clk),
    .D(net626),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7530_ (.CLK(clknet_leaf_5_clk),
    .D(net616),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7531_ (.CLK(clknet_leaf_10_clk),
    .D(net765),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7532_ (.CLK(clknet_leaf_77_clk),
    .D(net584),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7533_ (.CLK(clknet_leaf_78_clk),
    .D(net689),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7534_ (.CLK(clknet_leaf_12_clk),
    .D(net671),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7535_ (.CLK(clknet_leaf_45_clk),
    .D(net729),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7536_ (.CLK(clknet_leaf_11_clk),
    .D(net653),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7537_ (.CLK(clknet_leaf_13_clk),
    .D(net741),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7538_ (.CLK(clknet_leaf_46_clk),
    .D(net548),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7539_ (.CLK(clknet_leaf_19_clk),
    .D(net679),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7540_ (.CLK(clknet_leaf_27_clk),
    .D(net717),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7541_ (.CLK(clknet_leaf_48_clk),
    .D(net747),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7542_ (.CLK(clknet_leaf_66_clk),
    .D(net713),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7543_ (.CLK(clknet_leaf_61_clk),
    .D(net711),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7544_ (.CLK(clknet_leaf_67_clk),
    .D(net546),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7545_ (.CLK(clknet_leaf_66_clk),
    .D(net703),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7546_ (.CLK(clknet_leaf_48_clk),
    .D(net735),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7547_ (.CLK(clknet_leaf_62_clk),
    .D(net673),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7548_ (.CLK(clknet_leaf_61_clk),
    .D(net751),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7549_ (.CLK(clknet_leaf_55_clk),
    .D(net1514),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7550_ (.CLK(clknet_leaf_68_clk),
    .D(net622),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7551_ (.CLK(clknet_leaf_79_clk),
    .D(net731),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7552_ (.CLK(clknet_leaf_78_clk),
    .D(net767),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7553_ (.CLK(clknet_leaf_60_clk),
    .D(net737),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ));
 sky130_fd_sc_hd__dfxtp_2 _7554_ (.CLK(clknet_leaf_28_clk),
    .D(net2105),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7555_ (.CLK(clknet_leaf_35_clk),
    .D(net1178),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7556_ (.CLK(clknet_leaf_28_clk),
    .D(net2118),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7557_ (.CLK(clknet_leaf_28_clk),
    .D(net2145),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7558_ (.CLK(clknet_leaf_27_clk),
    .D(_0585_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ));
 sky130_fd_sc_hd__dfxtp_1 _7559_ (.CLK(clknet_leaf_24_clk),
    .D(net699),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _7560_ (.CLK(clknet_leaf_26_clk),
    .D(net556),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_2 _7561_ (.CLK(clknet_leaf_77_clk),
    .D(net677),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_2 _7562_ (.CLK(clknet_3_4_0_clk),
    .D(_0589_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_2 _7563_ (.CLK(clknet_leaf_54_clk),
    .D(_0590_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _7564_ (.CLK(clknet_leaf_82_clk),
    .D(_0591_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _7565_ (.CLK(clknet_3_0_0_clk),
    .D(_0592_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _7566_ (.CLK(clknet_leaf_26_clk),
    .D(_0593_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _7567_ (.CLK(clknet_leaf_25_clk),
    .D(_0594_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _7568_ (.CLK(clknet_leaf_12_clk),
    .D(_0595_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_2 _7569_ (.CLK(clknet_leaf_13_clk),
    .D(_0596_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_4 _7570_ (.CLK(clknet_leaf_38_clk),
    .D(_0597_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _7571_ (.CLK(clknet_leaf_78_clk),
    .D(_0598_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _7572_ (.CLK(clknet_leaf_13_clk),
    .D(_0599_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_2 _7573_ (.CLK(clknet_leaf_39_clk),
    .D(_0600_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_2 _7574_ (.CLK(clknet_leaf_79_clk),
    .D(_0601_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _7575_ (.CLK(clknet_leaf_5_clk),
    .D(_0602_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _7576_ (.CLK(clknet_leaf_61_clk),
    .D(_0603_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_2 _7577_ (.CLK(clknet_leaf_0_clk),
    .D(_0604_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_4 _7578_ (.CLK(clknet_leaf_4_clk),
    .D(_0605_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _7579_ (.CLK(clknet_3_4_0_clk),
    .D(_0606_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_4 _7580_ (.CLK(clknet_leaf_4_clk),
    .D(_0607_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _7581_ (.CLK(clknet_leaf_9_clk),
    .D(_0608_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _7582_ (.CLK(clknet_leaf_1_clk),
    .D(_0609_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _7583_ (.CLK(clknet_leaf_80_clk),
    .D(_0610_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _7584_ (.CLK(clknet_leaf_81_clk),
    .D(_0611_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _7585_ (.CLK(clknet_leaf_9_clk),
    .D(_0612_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _7586_ (.CLK(clknet_leaf_66_clk),
    .D(_0613_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _7587_ (.CLK(clknet_leaf_31_clk),
    .D(_0614_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _7588_ (.CLK(clknet_leaf_54_clk),
    .D(_0615_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _7589_ (.CLK(clknet_leaf_82_clk),
    .D(_0616_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _7590_ (.CLK(clknet_leaf_37_clk),
    .D(_0617_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _7591_ (.CLK(clknet_leaf_78_clk),
    .D(_0618_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _7592_ (.CLK(clknet_leaf_68_clk),
    .D(_0619_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _7593_ (.CLK(clknet_leaf_37_clk),
    .D(_0620_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _7594_ (.CLK(clknet_leaf_61_clk),
    .D(_0621_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _7595_ (.CLK(clknet_leaf_12_clk),
    .D(net723),
    .Q(\U_DATAPATH.U_EX_MEM.o_reg_write_M ));
 sky130_fd_sc_hd__dfxtp_1 _7596_ (.CLK(clknet_leaf_12_clk),
    .D(net1620),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7597_ (.CLK(clknet_leaf_12_clk),
    .D(net1283),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7598_ (.CLK(clknet_leaf_45_clk),
    .D(net2256),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_4 _7599_ (.CLK(clknet_leaf_46_clk),
    .D(_0626_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _7600_ (.CLK(clknet_leaf_45_clk),
    .D(net2339),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _7601_ (.CLK(clknet_leaf_16_clk),
    .D(_0628_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _7602_ (.CLK(clknet_leaf_16_clk),
    .D(_0629_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _7603_ (.CLK(clknet_leaf_22_clk),
    .D(_0630_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_4 _7604_ (.CLK(clknet_leaf_44_clk),
    .D(net2267),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _7605_ (.CLK(clknet_leaf_15_clk),
    .D(_0632_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_4 _7606_ (.CLK(clknet_leaf_3_clk),
    .D(_0633_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_4 _7607_ (.CLK(clknet_leaf_75_clk),
    .D(_0634_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _7608_ (.CLK(clknet_leaf_75_clk),
    .D(_0635_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _7609_ (.CLK(clknet_leaf_78_clk),
    .D(_0636_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_4 _7610_ (.CLK(clknet_leaf_75_clk),
    .D(_0637_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_4 _7611_ (.CLK(clknet_leaf_47_clk),
    .D(net2293),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_2 _7612_ (.CLK(clknet_leaf_11_clk),
    .D(_0639_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _7613_ (.CLK(clknet_leaf_15_clk),
    .D(net2326),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_4 _7614_ (.CLK(clknet_leaf_45_clk),
    .D(net2260),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_4 _7615_ (.CLK(clknet_leaf_47_clk),
    .D(net2295),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _7616_ (.CLK(clknet_leaf_19_clk),
    .D(_0643_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_4 _7617_ (.CLK(clknet_leaf_48_clk),
    .D(_0644_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_2 _7618_ (.CLK(clknet_leaf_48_clk),
    .D(_0645_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _7619_ (.CLK(clknet_leaf_72_clk),
    .D(_0646_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _7620_ (.CLK(clknet_leaf_73_clk),
    .D(_0647_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _7621_ (.CLK(clknet_leaf_73_clk),
    .D(_0648_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_4 _7622_ (.CLK(clknet_leaf_73_clk),
    .D(net2333),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _7623_ (.CLK(clknet_3_1_0_clk),
    .D(_0650_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_2 _7624_ (.CLK(clknet_leaf_70_clk),
    .D(_0651_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _7625_ (.CLK(clknet_leaf_48_clk),
    .D(_0652_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _7626_ (.CLK(clknet_leaf_76_clk),
    .D(_0653_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_4 _7627_ (.CLK(clknet_leaf_78_clk),
    .D(_0654_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_2 _7628_ (.CLK(clknet_leaf_75_clk),
    .D(_0655_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _7629_ (.CLK(clknet_leaf_48_clk),
    .D(net2299),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _7630_ (.CLK(clknet_leaf_20_clk),
    .D(net643),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7631_ (.CLK(clknet_leaf_11_clk),
    .D(net667),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7632_ (.CLK(clknet_leaf_10_clk),
    .D(net597),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7633_ (.CLK(clknet_leaf_11_clk),
    .D(net605),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7634_ (.CLK(clknet_leaf_44_clk),
    .D(net576),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7635_ (.CLK(clknet_leaf_15_clk),
    .D(net635),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7636_ (.CLK(clknet_leaf_5_clk),
    .D(net614),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7637_ (.CLK(clknet_leaf_10_clk),
    .D(net586),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7638_ (.CLK(clknet_leaf_0_clk),
    .D(net618),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7639_ (.CLK(clknet_leaf_78_clk),
    .D(net733),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7640_ (.CLK(clknet_leaf_12_clk),
    .D(net675),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7641_ (.CLK(clknet_leaf_45_clk),
    .D(net568),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7642_ (.CLK(clknet_leaf_11_clk),
    .D(net647),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7643_ (.CLK(clknet_leaf_13_clk),
    .D(net693),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7644_ (.CLK(clknet_leaf_17_clk),
    .D(net651),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7645_ (.CLK(clknet_leaf_19_clk),
    .D(net544),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7646_ (.CLK(clknet_leaf_27_clk),
    .D(net772),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7647_ (.CLK(clknet_leaf_48_clk),
    .D(net695),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7648_ (.CLK(clknet_leaf_66_clk),
    .D(net685),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7649_ (.CLK(clknet_leaf_61_clk),
    .D(net582),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7650_ (.CLK(clknet_leaf_68_clk),
    .D(net631),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7651_ (.CLK(clknet_leaf_66_clk),
    .D(net683),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7652_ (.CLK(clknet_leaf_48_clk),
    .D(net783),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7653_ (.CLK(clknet_leaf_62_clk),
    .D(net753),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7654_ (.CLK(clknet_leaf_61_clk),
    .D(net659),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7655_ (.CLK(clknet_leaf_61_clk),
    .D(net697),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7656_ (.CLK(clknet_leaf_68_clk),
    .D(net558),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7657_ (.CLK(clknet_leaf_79_clk),
    .D(net777),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7658_ (.CLK(clknet_leaf_78_clk),
    .D(net595),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7659_ (.CLK(clknet_leaf_61_clk),
    .D(net727),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7660_ (.CLK(clknet_leaf_28_clk),
    .D(_0687_),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7661_ (.CLK(clknet_leaf_20_clk),
    .D(_0688_),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7662_ (.CLK(clknet_leaf_27_clk),
    .D(net1309),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7663_ (.CLK(clknet_leaf_27_clk),
    .D(net1632),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7664_ (.CLK(clknet_leaf_35_clk),
    .D(net886),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7665_ (.CLK(clknet_leaf_36_clk),
    .D(net1064),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7666_ (.CLK(clknet_leaf_36_clk),
    .D(net908),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7667_ (.CLK(clknet_leaf_31_clk),
    .D(net980),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7668_ (.CLK(clknet_leaf_25_clk),
    .D(net1698),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7669_ (.CLK(clknet_leaf_24_clk),
    .D(net1267),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7670_ (.CLK(clknet_leaf_52_clk),
    .D(net1478),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7671_ (.CLK(clknet_leaf_41_clk),
    .D(net1330),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7672_ (.CLK(clknet_leaf_44_clk),
    .D(net1592),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7673_ (.CLK(clknet_leaf_30_clk),
    .D(net1273),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7674_ (.CLK(clknet_leaf_41_clk),
    .D(net1303),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7675_ (.CLK(clknet_leaf_69_clk),
    .D(net1673),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7676_ (.CLK(clknet_leaf_24_clk),
    .D(net1090),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7677_ (.CLK(clknet_leaf_54_clk),
    .D(net1414),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7678_ (.CLK(clknet_leaf_21_clk),
    .D(net1279),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7679_ (.CLK(clknet_leaf_21_clk),
    .D(net1516),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7680_ (.CLK(clknet_leaf_40_clk),
    .D(net1452),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7681_ (.CLK(clknet_leaf_20_clk),
    .D(net1628),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7682_ (.CLK(clknet_leaf_26_clk),
    .D(net1757),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7683_ (.CLK(clknet_leaf_48_clk),
    .D(net1317),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7684_ (.CLK(clknet_leaf_72_clk),
    .D(net1209),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7685_ (.CLK(clknet_leaf_55_clk),
    .D(net1522),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7686_ (.CLK(clknet_leaf_37_clk),
    .D(net1780),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7687_ (.CLK(clknet_leaf_63_clk),
    .D(net1000),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7688_ (.CLK(clknet_leaf_26_clk),
    .D(net1225),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7689_ (.CLK(clknet_leaf_64_clk),
    .D(net1374),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7690_ (.CLK(clknet_leaf_58_clk),
    .D(net1492),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7691_ (.CLK(clknet_leaf_39_clk),
    .D(net1056),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7692_ (.CLK(clknet_leaf_69_clk),
    .D(net994),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7693_ (.CLK(clknet_leaf_71_clk),
    .D(net1538),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7694_ (.CLK(clknet_leaf_49_clk),
    .D(net1376),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7695_ (.CLK(clknet_leaf_55_clk),
    .D(net1570),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7696_ (.CLK(clknet_leaf_34_clk),
    .D(net932),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7697_ (.CLK(clknet_leaf_33_clk),
    .D(net1344),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7698_ (.CLK(clknet_leaf_34_clk),
    .D(net1221),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7699_ (.CLK(clknet_leaf_34_clk),
    .D(net910),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7700_ (.CLK(clknet_leaf_27_clk),
    .D(net1751),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7701_ (.CLK(clknet_leaf_27_clk),
    .D(net1518),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7702_ (.CLK(clknet_leaf_52_clk),
    .D(net1366),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7703_ (.CLK(clknet_leaf_42_clk),
    .D(net1648),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7704_ (.CLK(clknet_leaf_44_clk),
    .D(net1358),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7705_ (.CLK(clknet_leaf_31_clk),
    .D(net968),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7706_ (.CLK(clknet_leaf_41_clk),
    .D(net1136),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7707_ (.CLK(clknet_leaf_71_clk),
    .D(net1338),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7708_ (.CLK(clknet_leaf_25_clk),
    .D(net1281),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7709_ (.CLK(clknet_leaf_54_clk),
    .D(net1410),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7710_ (.CLK(clknet_leaf_20_clk),
    .D(net1604),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7711_ (.CLK(clknet_leaf_19_clk),
    .D(net1086),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7712_ (.CLK(clknet_leaf_39_clk),
    .D(net1128),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7713_ (.CLK(clknet_leaf_43_clk),
    .D(net1418),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7714_ (.CLK(clknet_leaf_29_clk),
    .D(net1360),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7715_ (.CLK(clknet_leaf_50_clk),
    .D(net1520),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7716_ (.CLK(clknet_leaf_49_clk),
    .D(net1251),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7717_ (.CLK(clknet_leaf_54_clk),
    .D(net1116),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7718_ (.CLK(clknet_leaf_38_clk),
    .D(net1315),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7719_ (.CLK(clknet_leaf_58_clk),
    .D(net1444),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7720_ (.CLK(clknet_leaf_30_clk),
    .D(net1334),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7721_ (.CLK(clknet_leaf_64_clk),
    .D(net1510),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7722_ (.CLK(clknet_leaf_58_clk),
    .D(net1466),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7723_ (.CLK(clknet_leaf_52_clk),
    .D(net1370),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7724_ (.CLK(clknet_leaf_71_clk),
    .D(net1201),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7725_ (.CLK(clknet_leaf_64_clk),
    .D(net1915),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7726_ (.CLK(clknet_leaf_56_clk),
    .D(net1227),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7727_ (.CLK(clknet_leaf_55_clk),
    .D(net1687),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7728_ (.CLK(clknet_leaf_42_clk),
    .D(net775),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7729_ (.CLK(clknet_leaf_42_clk),
    .D(net829),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7730_ (.CLK(clknet_leaf_20_clk),
    .D(_0757_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7731_ (.CLK(clknet_leaf_11_clk),
    .D(_0758_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7732_ (.CLK(clknet_leaf_10_clk),
    .D(_0759_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7733_ (.CLK(clknet_leaf_11_clk),
    .D(_0760_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7734_ (.CLK(clknet_leaf_44_clk),
    .D(_0761_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7735_ (.CLK(clknet_leaf_15_clk),
    .D(_0762_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7736_ (.CLK(clknet_leaf_4_clk),
    .D(_0763_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7737_ (.CLK(clknet_leaf_10_clk),
    .D(_0764_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7738_ (.CLK(clknet_leaf_0_clk),
    .D(_0765_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7739_ (.CLK(clknet_leaf_78_clk),
    .D(_0766_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7740_ (.CLK(clknet_leaf_12_clk),
    .D(_0767_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7741_ (.CLK(clknet_leaf_15_clk),
    .D(_0768_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7742_ (.CLK(clknet_leaf_11_clk),
    .D(_0769_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7743_ (.CLK(clknet_leaf_13_clk),
    .D(_0770_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7744_ (.CLK(clknet_leaf_17_clk),
    .D(_0771_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7745_ (.CLK(clknet_leaf_19_clk),
    .D(_0772_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7746_ (.CLK(clknet_leaf_27_clk),
    .D(_0773_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7747_ (.CLK(clknet_leaf_48_clk),
    .D(_0774_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7748_ (.CLK(clknet_leaf_65_clk),
    .D(_0775_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7749_ (.CLK(clknet_leaf_62_clk),
    .D(_0776_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7750_ (.CLK(clknet_leaf_67_clk),
    .D(_0777_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7751_ (.CLK(clknet_leaf_67_clk),
    .D(_0778_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7752_ (.CLK(clknet_leaf_65_clk),
    .D(_0779_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7753_ (.CLK(clknet_leaf_62_clk),
    .D(_0780_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7754_ (.CLK(clknet_leaf_63_clk),
    .D(_0781_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7755_ (.CLK(clknet_leaf_61_clk),
    .D(_0782_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7756_ (.CLK(clknet_leaf_68_clk),
    .D(_0783_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7757_ (.CLK(clknet_leaf_79_clk),
    .D(_0784_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7758_ (.CLK(clknet_leaf_79_clk),
    .D(_0785_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7759_ (.CLK(clknet_leaf_61_clk),
    .D(_0786_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7760_ (.CLK(clknet_leaf_1_clk),
    .D(_0787_),
    .Q(\U_CONTROL_UNIT.i_jump_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7761_ (.CLK(clknet_leaf_1_clk),
    .D(_0788_),
    .Q(\U_CONTROL_UNIT.i_branch_EX ));
 sky130_fd_sc_hd__dfxtp_2 _7762_ (.CLK(clknet_leaf_4_clk),
    .D(_0789_),
    .Q(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7763_ (.CLK(clknet_leaf_12_clk),
    .D(_0790_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7764_ (.CLK(clknet_leaf_20_clk),
    .D(net1947),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7765_ (.CLK(clknet_leaf_20_clk),
    .D(_0792_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7766_ (.CLK(clknet_leaf_20_clk),
    .D(_0793_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7767_ (.CLK(clknet_leaf_35_clk),
    .D(_0794_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7768_ (.CLK(clknet_leaf_36_clk),
    .D(_0795_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7769_ (.CLK(clknet_leaf_42_clk),
    .D(_0796_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7770_ (.CLK(clknet_leaf_22_clk),
    .D(_0797_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7771_ (.CLK(clknet_leaf_23_clk),
    .D(_0798_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7772_ (.CLK(clknet_leaf_23_clk),
    .D(_0799_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7773_ (.CLK(clknet_leaf_41_clk),
    .D(_0800_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7774_ (.CLK(clknet_leaf_41_clk),
    .D(_0801_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7775_ (.CLK(clknet_leaf_44_clk),
    .D(_0802_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7776_ (.CLK(clknet_leaf_10_clk),
    .D(_0803_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7777_ (.CLK(clknet_leaf_47_clk),
    .D(_0804_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _7778_ (.CLK(clknet_leaf_70_clk),
    .D(_0805_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7779_ (.CLK(clknet_leaf_23_clk),
    .D(_0806_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7780_ (.CLK(clknet_leaf_51_clk),
    .D(_0807_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7781_ (.CLK(clknet_leaf_22_clk),
    .D(_0808_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7782_ (.CLK(clknet_leaf_17_clk),
    .D(_0809_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7783_ (.CLK(clknet_leaf_40_clk),
    .D(_0810_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7784_ (.CLK(clknet_leaf_43_clk),
    .D(_0811_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7785_ (.CLK(clknet_leaf_27_clk),
    .D(_0812_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7786_ (.CLK(clknet_leaf_47_clk),
    .D(_0813_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7787_ (.CLK(clknet_leaf_72_clk),
    .D(_0814_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7788_ (.CLK(clknet_leaf_56_clk),
    .D(_0815_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7789_ (.CLK(clknet_leaf_48_clk),
    .D(_0816_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7790_ (.CLK(clknet_leaf_64_clk),
    .D(_0817_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ));
 sky130_fd_sc_hd__dfxtp_4 _7791_ (.CLK(clknet_leaf_29_clk),
    .D(_0818_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7792_ (.CLK(clknet_leaf_63_clk),
    .D(_0819_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7793_ (.CLK(clknet_leaf_63_clk),
    .D(_0820_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7794_ (.CLK(clknet_leaf_50_clk),
    .D(_0821_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7795_ (.CLK(clknet_leaf_70_clk),
    .D(_0822_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7796_ (.CLK(clknet_leaf_69_clk),
    .D(_0823_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7797_ (.CLK(clknet_leaf_56_clk),
    .D(_0824_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7798_ (.CLK(clknet_leaf_56_clk),
    .D(_0825_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7799_ (.CLK(clknet_leaf_36_clk),
    .D(_0826_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7800_ (.CLK(clknet_leaf_36_clk),
    .D(_0827_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7801_ (.CLK(clknet_leaf_42_clk),
    .D(_0828_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7802_ (.CLK(clknet_leaf_22_clk),
    .D(_0829_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7803_ (.CLK(clknet_leaf_23_clk),
    .D(_0830_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7804_ (.CLK(clknet_leaf_23_clk),
    .D(_0831_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7805_ (.CLK(clknet_leaf_41_clk),
    .D(_0832_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7806_ (.CLK(clknet_leaf_42_clk),
    .D(_0833_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7807_ (.CLK(clknet_leaf_45_clk),
    .D(_0834_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7808_ (.CLK(clknet_leaf_23_clk),
    .D(_0835_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7809_ (.CLK(clknet_leaf_47_clk),
    .D(_0836_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7810_ (.CLK(clknet_leaf_70_clk),
    .D(_0837_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7811_ (.CLK(clknet_leaf_23_clk),
    .D(_0838_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7812_ (.CLK(clknet_leaf_51_clk),
    .D(_0839_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7813_ (.CLK(clknet_leaf_22_clk),
    .D(_0840_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7814_ (.CLK(clknet_leaf_14_clk),
    .D(_0841_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7815_ (.CLK(clknet_leaf_40_clk),
    .D(_0842_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7816_ (.CLK(clknet_leaf_43_clk),
    .D(_0843_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7817_ (.CLK(clknet_leaf_27_clk),
    .D(_0844_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7818_ (.CLK(clknet_leaf_47_clk),
    .D(_0845_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7819_ (.CLK(clknet_leaf_64_clk),
    .D(_0846_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7820_ (.CLK(clknet_leaf_56_clk),
    .D(_0847_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7821_ (.CLK(clknet_leaf_36_clk),
    .D(_0848_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7822_ (.CLK(clknet_leaf_64_clk),
    .D(_0849_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7823_ (.CLK(clknet_leaf_29_clk),
    .D(_0850_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7824_ (.CLK(clknet_leaf_49_clk),
    .D(_0851_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7825_ (.CLK(clknet_leaf_64_clk),
    .D(_0852_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7826_ (.CLK(clknet_leaf_51_clk),
    .D(_0853_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7827_ (.CLK(clknet_leaf_78_clk),
    .D(_0854_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7828_ (.CLK(clknet_leaf_70_clk),
    .D(_0855_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7829_ (.CLK(clknet_leaf_48_clk),
    .D(_0856_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7830_ (.CLK(clknet_leaf_56_clk),
    .D(_0857_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7831_ (.CLK(clknet_leaf_28_clk),
    .D(_0858_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7832_ (.CLK(clknet_leaf_28_clk),
    .D(_0859_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7833_ (.CLK(clknet_leaf_28_clk),
    .D(_0860_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7834_ (.CLK(clknet_leaf_28_clk),
    .D(_0861_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7835_ (.CLK(clknet_leaf_27_clk),
    .D(_0862_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7836_ (.CLK(clknet_leaf_27_clk),
    .D(_0863_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7837_ (.CLK(clknet_leaf_27_clk),
    .D(_0864_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7838_ (.CLK(clknet_leaf_28_clk),
    .D(_0865_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7839_ (.CLK(clknet_leaf_44_clk),
    .D(net823),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7840_ (.CLK(clknet_leaf_22_clk),
    .D(net770),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7841_ (.CLK(clknet_leaf_18_clk),
    .D(net850),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7842_ (.CLK(clknet_leaf_11_clk),
    .D(net813),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7843_ (.CLK(clknet_leaf_41_clk),
    .D(net842),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7844_ (.CLK(clknet_leaf_4_clk),
    .D(net797),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7845_ (.CLK(clknet_leaf_4_clk),
    .D(net866),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7846_ (.CLK(clknet_leaf_10_clk),
    .D(net805),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7847_ (.CLK(clknet_leaf_2_clk),
    .D(net1011),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7848_ (.CLK(clknet_leaf_13_clk),
    .D(net888),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7849_ (.CLK(clknet_leaf_12_clk),
    .D(net844),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7850_ (.CLK(clknet_leaf_42_clk),
    .D(net562),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7851_ (.CLK(clknet_leaf_10_clk),
    .D(net833),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7852_ (.CLK(clknet_leaf_14_clk),
    .D(net572),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7853_ (.CLK(clknet_leaf_19_clk),
    .D(net542),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7854_ (.CLK(clknet_leaf_43_clk),
    .D(net792),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7855_ (.CLK(clknet_leaf_23_clk),
    .D(net610),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7856_ (.CLK(clknet_leaf_47_clk),
    .D(net836),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7857_ (.CLK(clknet_leaf_66_clk),
    .D(net892),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7858_ (.CLK(clknet_leaf_62_clk),
    .D(net870),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7859_ (.CLK(clknet_leaf_67_clk),
    .D(net846),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7860_ (.CLK(clknet_leaf_67_clk),
    .D(net898),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7861_ (.CLK(clknet_leaf_65_clk),
    .D(net975),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7862_ (.CLK(clknet_leaf_61_clk),
    .D(net817),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7863_ (.CLK(clknet_leaf_61_clk),
    .D(net884),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7864_ (.CLK(clknet_leaf_69_clk),
    .D(net645),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7865_ (.CLK(clknet_leaf_68_clk),
    .D(net880),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7866_ (.CLK(clknet_leaf_79_clk),
    .D(net564),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7867_ (.CLK(clknet_leaf_79_clk),
    .D(net801),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7868_ (.CLK(clknet_leaf_63_clk),
    .D(net819),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7869_ (.CLK(clknet_leaf_20_clk),
    .D(net874),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7870_ (.CLK(clknet_leaf_11_clk),
    .D(net840),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7871_ (.CLK(clknet_leaf_12_clk),
    .D(net629),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7872_ (.CLK(clknet_leaf_12_clk),
    .D(net607),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7873_ (.CLK(clknet_leaf_19_clk),
    .D(net552),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7874_ (.CLK(clknet_leaf_13_clk),
    .D(net876),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7875_ (.CLK(clknet_leaf_5_clk),
    .D(net779),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7876_ (.CLK(clknet_leaf_12_clk),
    .D(net815),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7877_ (.CLK(clknet_leaf_0_clk),
    .D(net755),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7878_ (.CLK(clknet_leaf_78_clk),
    .D(net540),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7879_ (.CLK(clknet_leaf_12_clk),
    .D(net831),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7880_ (.CLK(clknet_leaf_14_clk),
    .D(net560),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7881_ (.CLK(clknet_leaf_11_clk),
    .D(net848),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7882_ (.CLK(clknet_leaf_13_clk),
    .D(net857),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7883_ (.CLK(clknet_leaf_17_clk),
    .D(net803),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7884_ (.CLK(clknet_leaf_18_clk),
    .D(net794),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7885_ (.CLK(clknet_leaf_27_clk),
    .D(net759),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7886_ (.CLK(clknet_leaf_48_clk),
    .D(net719),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7887_ (.CLK(clknet_leaf_66_clk),
    .D(net811),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7888_ (.CLK(clknet_leaf_62_clk),
    .D(net657),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7889_ (.CLK(clknet_leaf_68_clk),
    .D(net864),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7890_ (.CLK(clknet_leaf_66_clk),
    .D(net862),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7891_ (.CLK(clknet_leaf_48_clk),
    .D(_0918_),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7892_ (.CLK(clknet_leaf_62_clk),
    .D(net825),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7893_ (.CLK(clknet_leaf_61_clk),
    .D(net859),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7894_ (.CLK(clknet_leaf_61_clk),
    .D(net612),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7895_ (.CLK(clknet_leaf_80_clk),
    .D(net743),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7896_ (.CLK(clknet_leaf_79_clk),
    .D(net838),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7897_ (.CLK(clknet_leaf_79_clk),
    .D(net799),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7898_ (.CLK(clknet_leaf_61_clk),
    .D(net566),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7899_ (.CLK(clknet_leaf_12_clk),
    .D(_0926_),
    .Q(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7900_ (.CLK(clknet_leaf_12_clk),
    .D(_0927_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7901_ (.CLK(clknet_leaf_4_clk),
    .D(_0928_),
    .Q(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7902_ (.CLK(clknet_leaf_2_clk),
    .D(_0929_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ));
 sky130_fd_sc_hd__dfxtp_4 _7903_ (.CLK(clknet_leaf_4_clk),
    .D(_0930_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7904_ (.CLK(clknet_leaf_33_clk),
    .D(net1170),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7905_ (.CLK(clknet_leaf_33_clk),
    .D(net1352),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7906_ (.CLK(clknet_leaf_34_clk),
    .D(net1048),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7907_ (.CLK(clknet_leaf_34_clk),
    .D(net1033),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7908_ (.CLK(clknet_leaf_27_clk),
    .D(net1476),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7909_ (.CLK(clknet_leaf_27_clk),
    .D(net1428),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7910_ (.CLK(clknet_leaf_52_clk),
    .D(net1326),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7911_ (.CLK(clknet_leaf_42_clk),
    .D(net1420),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7912_ (.CLK(clknet_leaf_41_clk),
    .D(net1380),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7913_ (.CLK(clknet_leaf_32_clk),
    .D(net1036),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7914_ (.CLK(clknet_leaf_51_clk),
    .D(net1726),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7915_ (.CLK(clknet_leaf_72_clk),
    .D(net1237),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7916_ (.CLK(clknet_leaf_23_clk),
    .D(net1679),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7917_ (.CLK(clknet_leaf_54_clk),
    .D(net1263),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7918_ (.CLK(clknet_leaf_21_clk),
    .D(net1564),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7919_ (.CLK(clknet_leaf_19_clk),
    .D(net1245),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7920_ (.CLK(clknet_leaf_40_clk),
    .D(net1743),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7921_ (.CLK(clknet_leaf_42_clk),
    .D(net1829),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7922_ (.CLK(clknet_leaf_26_clk),
    .D(net1661),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7923_ (.CLK(clknet_leaf_51_clk),
    .D(net1802),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7924_ (.CLK(clknet_leaf_49_clk),
    .D(net1054),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7925_ (.CLK(clknet_leaf_55_clk),
    .D(net1663),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7926_ (.CLK(clknet_leaf_37_clk),
    .D(net1454),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7927_ (.CLK(clknet_leaf_57_clk),
    .D(net1142),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7928_ (.CLK(clknet_leaf_29_clk),
    .D(net1618),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7929_ (.CLK(clknet_leaf_57_clk),
    .D(net1154),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7930_ (.CLK(clknet_leaf_59_clk),
    .D(net1480),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7931_ (.CLK(clknet_leaf_40_clk),
    .D(net1546),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7932_ (.CLK(clknet_leaf_71_clk),
    .D(net1512),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7933_ (.CLK(clknet_leaf_64_clk),
    .D(net1640),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7934_ (.CLK(clknet_leaf_56_clk),
    .D(net1887),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7935_ (.CLK(clknet_leaf_55_clk),
    .D(net1426),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7936_ (.CLK(clknet_leaf_34_clk),
    .D(net912),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7937_ (.CLK(clknet_leaf_34_clk),
    .D(net940),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7938_ (.CLK(clknet_leaf_34_clk),
    .D(net853),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7939_ (.CLK(clknet_leaf_29_clk),
    .D(net936),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7940_ (.CLK(clknet_leaf_27_clk),
    .D(net1689),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7941_ (.CLK(clknet_leaf_21_clk),
    .D(net1382),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7942_ (.CLK(clknet_leaf_51_clk),
    .D(net1616),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7943_ (.CLK(clknet_leaf_42_clk),
    .D(net1724),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7944_ (.CLK(clknet_leaf_44_clk),
    .D(net1213),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7945_ (.CLK(clknet_leaf_29_clk),
    .D(net1269),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7946_ (.CLK(clknet_leaf_47_clk),
    .D(net1602),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7947_ (.CLK(clknet_leaf_70_clk),
    .D(net1524),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7948_ (.CLK(clknet_leaf_23_clk),
    .D(net1490),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7949_ (.CLK(clknet_leaf_50_clk),
    .D(net1060),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7950_ (.CLK(clknet_leaf_21_clk),
    .D(net1199),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7951_ (.CLK(clknet_leaf_18_clk),
    .D(net992),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7952_ (.CLK(clknet_leaf_40_clk),
    .D(net1422),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7953_ (.CLK(clknet_leaf_43_clk),
    .D(net1172),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7954_ (.CLK(clknet_leaf_26_clk),
    .D(net1691),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7955_ (.CLK(clknet_leaf_51_clk),
    .D(net1634),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7956_ (.CLK(clknet_leaf_48_clk),
    .D(net1582),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7957_ (.CLK(clknet_leaf_56_clk),
    .D(net1346),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7958_ (.CLK(clknet_leaf_42_clk),
    .D(net1657),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7959_ (.CLK(clknet_leaf_57_clk),
    .D(net1293),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7960_ (.CLK(clknet_leaf_29_clk),
    .D(net1176),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7961_ (.CLK(clknet_leaf_57_clk),
    .D(net1277),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7962_ (.CLK(clknet_leaf_57_clk),
    .D(net1287),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7963_ (.CLK(clknet_leaf_41_clk),
    .D(net1207),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7964_ (.CLK(clknet_leaf_70_clk),
    .D(net1540),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7965_ (.CLK(clknet_leaf_71_clk),
    .D(net1416),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7966_ (.CLK(clknet_leaf_56_clk),
    .D(net1532),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7967_ (.CLK(clknet_leaf_56_clk),
    .D(net1390),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7968_ (.CLK(clknet_leaf_34_clk),
    .D(net1094),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7969_ (.CLK(clknet_leaf_34_clk),
    .D(net960),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7970_ (.CLK(clknet_leaf_34_clk),
    .D(net902),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7971_ (.CLK(clknet_leaf_29_clk),
    .D(net948),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7972_ (.CLK(clknet_leaf_27_clk),
    .D(net1328),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7973_ (.CLK(clknet_leaf_23_clk),
    .D(net1796),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7974_ (.CLK(clknet_leaf_51_clk),
    .D(net1586),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7975_ (.CLK(clknet_leaf_42_clk),
    .D(net1368),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7976_ (.CLK(clknet_leaf_44_clk),
    .D(net1124),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7977_ (.CLK(clknet_leaf_29_clk),
    .D(net1249),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7978_ (.CLK(clknet_leaf_47_clk),
    .D(net1438),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7979_ (.CLK(clknet_leaf_70_clk),
    .D(net1636),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7980_ (.CLK(clknet_leaf_23_clk),
    .D(net1392),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7981_ (.CLK(clknet_leaf_52_clk),
    .D(net1626),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7982_ (.CLK(clknet_leaf_21_clk),
    .D(net1253),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7983_ (.CLK(clknet_leaf_18_clk),
    .D(net1229),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7984_ (.CLK(clknet_leaf_40_clk),
    .D(net1470),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7985_ (.CLK(clknet_leaf_43_clk),
    .D(net1009),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7986_ (.CLK(clknet_leaf_27_clk),
    .D(net1482),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7987_ (.CLK(clknet_leaf_51_clk),
    .D(net1464),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7988_ (.CLK(clknet_leaf_72_clk),
    .D(net1456),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7989_ (.CLK(clknet_leaf_56_clk),
    .D(net1782),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7990_ (.CLK(clknet_leaf_42_clk),
    .D(net1736),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7991_ (.CLK(clknet_leaf_57_clk),
    .D(net1235),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7992_ (.CLK(clknet_leaf_29_clk),
    .D(net1695),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7993_ (.CLK(clknet_leaf_64_clk),
    .D(net1502),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7994_ (.CLK(clknet_leaf_57_clk),
    .D(net1430),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7995_ (.CLK(clknet_leaf_41_clk),
    .D(net1243),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7996_ (.CLK(clknet_leaf_70_clk),
    .D(net1574),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7997_ (.CLK(clknet_leaf_71_clk),
    .D(net1450),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7998_ (.CLK(clknet_leaf_56_clk),
    .D(net1265),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7999_ (.CLK(clknet_leaf_56_clk),
    .D(net1486),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8000_ (.CLK(net505),
    .D(_0000_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8001_ (.CLK(net506),
    .D(_0011_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8002_ (.CLK(net507),
    .D(_0022_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8003_ (.CLK(net508),
    .D(_0025_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8004_ (.CLK(net509),
    .D(_0026_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8005_ (.CLK(net510),
    .D(_0027_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8006_ (.CLK(net511),
    .D(_0028_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8007_ (.CLK(net512),
    .D(_0029_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8008_ (.CLK(net513),
    .D(_0030_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8009_ (.CLK(net514),
    .D(_0031_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8010_ (.CLK(net515),
    .D(_0001_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8011_ (.CLK(net516),
    .D(_0002_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8012_ (.CLK(net517),
    .D(_0003_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8013_ (.CLK(net518),
    .D(_0004_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8014_ (.CLK(net519),
    .D(_0005_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8015_ (.CLK(net520),
    .D(_0006_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8016_ (.CLK(net521),
    .D(_0007_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8017_ (.CLK(net522),
    .D(_0008_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8018_ (.CLK(net523),
    .D(_0009_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(net524),
    .D(_0010_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8020_ (.CLK(net525),
    .D(_0012_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(net526),
    .D(_0013_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8022_ (.CLK(net527),
    .D(_0014_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(net528),
    .D(_0015_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8024_ (.CLK(net529),
    .D(_0016_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(net530),
    .D(_0017_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(net531),
    .D(_0018_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(net532),
    .D(_0019_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(net533),
    .D(_0020_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8029_ (.CLK(net534),
    .D(_0021_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(net535),
    .D(_0023_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8031_ (.CLK(net536),
    .D(_0024_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(clknet_leaf_35_clk),
    .D(net894),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(clknet_leaf_36_clk),
    .D(net1700),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(clknet_leaf_35_clk),
    .D(net926),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(clknet_leaf_32_clk),
    .D(net1566),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(clknet_leaf_25_clk),
    .D(net1092),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(clknet_leaf_24_clk),
    .D(net1070),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(clknet_leaf_53_clk),
    .D(net1568),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(clknet_leaf_41_clk),
    .D(net1130),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(clknet_leaf_45_clk),
    .D(net1412),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(clknet_leaf_31_clk),
    .D(net966),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(clknet_leaf_41_clk),
    .D(net1174),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(clknet_leaf_69_clk),
    .D(net1548),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8044_ (.CLK(clknet_leaf_24_clk),
    .D(net1023),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8045_ (.CLK(clknet_leaf_54_clk),
    .D(net1323),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(clknet_leaf_21_clk),
    .D(net1112),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(clknet_leaf_21_clk),
    .D(net1458),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(clknet_leaf_39_clk),
    .D(net1160),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(clknet_leaf_20_clk),
    .D(net1295),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8050_ (.CLK(clknet_leaf_26_clk),
    .D(net1594),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8051_ (.CLK(clknet_leaf_50_clk),
    .D(net1186),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8052_ (.CLK(clknet_leaf_49_clk),
    .D(net1066),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8053_ (.CLK(clknet_leaf_54_clk),
    .D(net1180),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8054_ (.CLK(clknet_leaf_37_clk),
    .D(net1082),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8055_ (.CLK(clknet_leaf_58_clk),
    .D(net1100),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8056_ (.CLK(clknet_leaf_29_clk),
    .D(net1534),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8057_ (.CLK(clknet_leaf_64_clk),
    .D(net1710),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8058_ (.CLK(clknet_leaf_60_clk),
    .D(net1062),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8059_ (.CLK(clknet_leaf_39_clk),
    .D(net1021),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8060_ (.CLK(clknet_leaf_70_clk),
    .D(net1215),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8061_ (.CLK(clknet_leaf_65_clk),
    .D(net946),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8062_ (.CLK(clknet_leaf_49_clk),
    .D(net998),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8063_ (.CLK(clknet_leaf_55_clk),
    .D(net1572),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8064_ (.CLK(clknet_leaf_33_clk),
    .D(net1080),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8065_ (.CLK(clknet_leaf_37_clk),
    .D(net1006),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(clknet_leaf_36_clk),
    .D(net1588),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8067_ (.CLK(clknet_leaf_32_clk),
    .D(net1432),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8068_ (.CLK(clknet_leaf_25_clk),
    .D(net1498),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8069_ (.CLK(clknet_leaf_24_clk),
    .D(net1526),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8070_ (.CLK(clknet_leaf_53_clk),
    .D(net1291),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8071_ (.CLK(clknet_leaf_40_clk),
    .D(net1193),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8072_ (.CLK(clknet_leaf_45_clk),
    .D(net1530),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8073_ (.CLK(clknet_leaf_30_clk),
    .D(net1554),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8074_ (.CLK(clknet_leaf_51_clk),
    .D(net1638),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8075_ (.CLK(clknet_leaf_69_clk),
    .D(net1550),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8076_ (.CLK(clknet_leaf_23_clk),
    .D(net1528),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8077_ (.CLK(clknet_leaf_53_clk),
    .D(net1239),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8078_ (.CLK(clknet_leaf_21_clk),
    .D(net1600),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8079_ (.CLK(clknet_leaf_18_clk),
    .D(net1152),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8080_ (.CLK(clknet_leaf_39_clk),
    .D(net1025),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8081_ (.CLK(clknet_leaf_20_clk),
    .D(net1622),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(clknet_leaf_26_clk),
    .D(net1749),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8083_ (.CLK(clknet_leaf_51_clk),
    .D(net1794),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8084_ (.CLK(clknet_leaf_57_clk),
    .D(net1402),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8085_ (.CLK(clknet_leaf_55_clk),
    .D(net1677),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8086_ (.CLK(clknet_leaf_38_clk),
    .D(net1440),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8087_ (.CLK(clknet_leaf_60_clk),
    .D(net1078),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8088_ (.CLK(clknet_leaf_30_clk),
    .D(net1650),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8089_ (.CLK(clknet_leaf_63_clk),
    .D(net1255),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8090_ (.CLK(clknet_leaf_60_clk),
    .D(net1074),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8091_ (.CLK(clknet_leaf_53_clk),
    .D(net1400),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8092_ (.CLK(clknet_leaf_69_clk),
    .D(net1027),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8093_ (.CLK(clknet_leaf_64_clk),
    .D(net1386),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8094_ (.CLK(clknet_leaf_50_clk),
    .D(net1448),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8095_ (.CLK(clknet_leaf_59_clk),
    .D(net1722),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8096_ (.CLK(clknet_leaf_36_clk),
    .D(net1311),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8097_ (.CLK(clknet_leaf_36_clk),
    .D(net996),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8098_ (.CLK(clknet_leaf_35_clk),
    .D(net872),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8099_ (.CLK(clknet_leaf_31_clk),
    .D(net988),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8100_ (.CLK(clknet_leaf_24_clk),
    .D(net1257),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8101_ (.CLK(clknet_leaf_24_clk),
    .D(net1140),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8102_ (.CLK(clknet_leaf_52_clk),
    .D(net1624),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8103_ (.CLK(clknet_leaf_41_clk),
    .D(net1231),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8104_ (.CLK(clknet_leaf_45_clk),
    .D(net1203),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8105_ (.CLK(clknet_leaf_30_clk),
    .D(net1096),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8106_ (.CLK(clknet_leaf_41_clk),
    .D(net1205),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8107_ (.CLK(clknet_leaf_69_clk),
    .D(net1148),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8108_ (.CLK(clknet_leaf_23_clk),
    .D(net1562),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8109_ (.CLK(clknet_leaf_54_clk),
    .D(net1197),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8110_ (.CLK(clknet_leaf_21_clk),
    .D(net1068),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8111_ (.CLK(clknet_leaf_22_clk),
    .D(net1275),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8112_ (.CLK(clknet_leaf_39_clk),
    .D(net1013),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8113_ (.CLK(clknet_leaf_20_clk),
    .D(net1610),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8114_ (.CLK(clknet_leaf_25_clk),
    .D(net1321),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8115_ (.CLK(clknet_leaf_48_clk),
    .D(net1642),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8116_ (.CLK(clknet_leaf_72_clk),
    .D(net1158),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8117_ (.CLK(clknet_leaf_54_clk),
    .D(net1211),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8118_ (.CLK(clknet_leaf_37_clk),
    .D(net1076),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8119_ (.CLK(clknet_leaf_58_clk),
    .D(net1552),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8120_ (.CLK(clknet_leaf_26_clk),
    .D(net1340),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8121_ (.CLK(clknet_leaf_64_clk),
    .D(net1703),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8122_ (.CLK(clknet_leaf_58_clk),
    .D(net1590),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8123_ (.CLK(clknet_leaf_39_clk),
    .D(net1004),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8124_ (.CLK(clknet_leaf_69_clk),
    .D(net1342),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8125_ (.CLK(clknet_leaf_71_clk),
    .D(net1110),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8126_ (.CLK(clknet_leaf_49_clk),
    .D(net1434),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8127_ (.CLK(clknet_leaf_58_clk),
    .D(net1108),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8128_ (.CLK(clknet_leaf_34_clk),
    .D(net918),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8129_ (.CLK(clknet_leaf_36_clk),
    .D(net1285),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8130_ (.CLK(clknet_leaf_34_clk),
    .D(net1424),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8131_ (.CLK(clknet_leaf_29_clk),
    .D(net868),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8132_ (.CLK(clknet_leaf_26_clk),
    .D(net1734),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8133_ (.CLK(clknet_leaf_21_clk),
    .D(net1104),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8134_ (.CLK(clknet_leaf_52_clk),
    .D(net1120),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8135_ (.CLK(clknet_leaf_42_clk),
    .D(net1446),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8136_ (.CLK(clknet_leaf_41_clk),
    .D(net1496),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8137_ (.CLK(clknet_leaf_31_clk),
    .D(net1046),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8138_ (.CLK(clknet_leaf_51_clk),
    .D(net1708),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8139_ (.CLK(clknet_leaf_73_clk),
    .D(net928),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8140_ (.CLK(clknet_leaf_23_clk),
    .D(net1867),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8141_ (.CLK(clknet_leaf_51_clk),
    .D(net1404),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8142_ (.CLK(clknet_leaf_21_clk),
    .D(net1560),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8143_ (.CLK(clknet_leaf_18_clk),
    .D(net1031),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8144_ (.CLK(clknet_leaf_40_clk),
    .D(net1378),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8145_ (.CLK(clknet_leaf_42_clk),
    .D(net1598),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8146_ (.CLK(clknet_leaf_26_clk),
    .D(net1713),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8147_ (.CLK(clknet_leaf_50_clk),
    .D(net1348),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8148_ (.CLK(clknet_leaf_48_clk),
    .D(net1188),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8149_ (.CLK(clknet_leaf_55_clk),
    .D(net1408),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8150_ (.CLK(clknet_leaf_38_clk),
    .D(net1394),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8151_ (.CLK(clknet_leaf_57_clk),
    .D(net952),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8152_ (.CLK(clknet_leaf_29_clk),
    .D(net1659),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8153_ (.CLK(clknet_leaf_57_clk),
    .D(net1233),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8154_ (.CLK(clknet_leaf_59_clk),
    .D(net1017),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8155_ (.CLK(clknet_leaf_40_clk),
    .D(net1608),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8156_ (.CLK(clknet_leaf_70_clk),
    .D(net1504),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8157_ (.CLK(clknet_leaf_72_clk),
    .D(net1442),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8158_ (.CLK(clknet_leaf_56_clk),
    .D(net1106),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8159_ (.CLK(clknet_leaf_55_clk),
    .D(net1362),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8160_ (.CLK(clknet_leaf_44_clk),
    .D(net977),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8161_ (.CLK(clknet_leaf_22_clk),
    .D(net904),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8162_ (.CLK(clknet_leaf_18_clk),
    .D(net757),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8163_ (.CLK(clknet_leaf_11_clk),
    .D(net821),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8164_ (.CLK(clknet_leaf_41_clk),
    .D(net788),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8165_ (.CLK(clknet_leaf_4_clk),
    .D(net942),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8166_ (.CLK(clknet_leaf_4_clk),
    .D(net954),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8167_ (.CLK(clknet_leaf_10_clk),
    .D(net964),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8168_ (.CLK(clknet_leaf_2_clk),
    .D(net807),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8169_ (.CLK(clknet_leaf_13_clk),
    .D(net1102),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8170_ (.CLK(clknet_leaf_12_clk),
    .D(net990),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8171_ (.CLK(clknet_leaf_43_clk),
    .D(net906),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8172_ (.CLK(clknet_leaf_10_clk),
    .D(net1002),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8173_ (.CLK(clknet_leaf_13_clk),
    .D(net1084),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8174_ (.CLK(clknet_leaf_17_clk),
    .D(net916),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8175_ (.CLK(clknet_leaf_43_clk),
    .D(net938),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8176_ (.CLK(clknet_leaf_10_clk),
    .D(net982),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8177_ (.CLK(clknet_leaf_47_clk),
    .D(net1144),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8178_ (.CLK(clknet_leaf_66_clk),
    .D(net956),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8179_ (.CLK(clknet_leaf_62_clk),
    .D(net973),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8180_ (.CLK(clknet_leaf_67_clk),
    .D(net944),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8181_ (.CLK(clknet_leaf_67_clk),
    .D(net924),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8182_ (.CLK(clknet_leaf_66_clk),
    .D(net1044),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8183_ (.CLK(clknet_leaf_61_clk),
    .D(net669),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8184_ (.CLK(clknet_leaf_61_clk),
    .D(net1019),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8185_ (.CLK(clknet_leaf_68_clk),
    .D(net930),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8186_ (.CLK(clknet_leaf_68_clk),
    .D(net914),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8187_ (.CLK(clknet_leaf_80_clk),
    .D(net855),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8188_ (.CLK(clknet_leaf_79_clk),
    .D(net934),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8189_ (.CLK(clknet_leaf_63_clk),
    .D(net900),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ));
 sky130_fd_sc_hd__dfxtp_2 _8190_ (.CLK(clknet_leaf_78_clk),
    .D(_1185_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8191_ (.CLK(clknet_leaf_4_clk),
    .D(_1186_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8192_ (.CLK(clknet_leaf_4_clk),
    .D(_1187_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8193_ (.CLK(clknet_leaf_4_clk),
    .D(_1188_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8194_ (.CLK(clknet_leaf_4_clk),
    .D(_1189_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8195_ (.CLK(clknet_leaf_8_clk),
    .D(_1190_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8196_ (.CLK(clknet_leaf_4_clk),
    .D(_1191_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(clknet_leaf_32_clk),
    .D(_1192_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(clknet_leaf_8_clk),
    .D(_1193_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8199_ (.CLK(clknet_leaf_1_clk),
    .D(_1194_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ));
 sky130_fd_sc_hd__dfxtp_2 _8200_ (.CLK(clknet_leaf_79_clk),
    .D(_1195_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8201_ (.CLK(clknet_leaf_4_clk),
    .D(_1196_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(clknet_leaf_3_clk),
    .D(_1197_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8203_ (.CLK(clknet_leaf_9_clk),
    .D(_1198_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(clknet_leaf_54_clk),
    .D(_1199_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_4 _8205_ (.CLK(clknet_leaf_66_clk),
    .D(_1200_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8206_ (.CLK(clknet_leaf_68_clk),
    .D(_1201_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8207_ (.CLK(clknet_leaf_37_clk),
    .D(_1202_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(clknet_leaf_32_clk),
    .D(_1203_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8209_ (.CLK(clknet_leaf_55_clk),
    .D(_1204_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8210_ (.CLK(clknet_leaf_32_clk),
    .D(_1205_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8211_ (.CLK(clknet_leaf_59_clk),
    .D(_1206_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(clknet_leaf_37_clk),
    .D(_1207_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8213_ (.CLK(clknet_leaf_0_clk),
    .D(_1208_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8214_ (.CLK(clknet_leaf_67_clk),
    .D(_1209_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(clknet_leaf_37_clk),
    .D(_1210_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8216_ (.CLK(clknet_leaf_81_clk),
    .D(_1211_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(clknet_leaf_10_clk),
    .D(_1212_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ));
 sky130_fd_sc_hd__dfxtp_4 _8218_ (.CLK(clknet_leaf_61_clk),
    .D(_1213_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(clknet_leaf_2_clk),
    .D(_1214_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(clknet_leaf_20_clk),
    .D(_1215_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(clknet_leaf_11_clk),
    .D(_1216_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(clknet_leaf_10_clk),
    .D(_1217_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(clknet_leaf_11_clk),
    .D(_1218_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(clknet_leaf_14_clk),
    .D(_1219_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(clknet_leaf_13_clk),
    .D(net950),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8226_ (.CLK(clknet_leaf_5_clk),
    .D(_1221_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(clknet_leaf_12_clk),
    .D(_1222_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(clknet_leaf_0_clk),
    .D(net2044),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(clknet_leaf_77_clk),
    .D(_1224_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8230_ (.CLK(clknet_leaf_12_clk),
    .D(_1225_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8231_ (.CLK(clknet_leaf_15_clk),
    .D(_1226_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(clknet_leaf_11_clk),
    .D(_1227_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(clknet_leaf_13_clk),
    .D(_1228_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(clknet_leaf_17_clk),
    .D(_1229_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8235_ (.CLK(clknet_leaf_18_clk),
    .D(_1230_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8236_ (.CLK(clknet_leaf_21_clk),
    .D(net890),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8237_ (.CLK(clknet_leaf_47_clk),
    .D(_1232_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8238_ (.CLK(clknet_leaf_66_clk),
    .D(_1233_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8239_ (.CLK(clknet_leaf_66_clk),
    .D(_1234_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8240_ (.CLK(clknet_leaf_67_clk),
    .D(_1235_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8241_ (.CLK(clknet_leaf_66_clk),
    .D(_1236_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8242_ (.CLK(clknet_leaf_66_clk),
    .D(_1237_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8243_ (.CLK(clknet_leaf_62_clk),
    .D(_1238_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8244_ (.CLK(clknet_leaf_61_clk),
    .D(net1956),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8245_ (.CLK(clknet_leaf_62_clk),
    .D(_1240_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8246_ (.CLK(clknet_leaf_80_clk),
    .D(net2026),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8247_ (.CLK(clknet_leaf_79_clk),
    .D(_1242_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8248_ (.CLK(clknet_leaf_79_clk),
    .D(_1243_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8249_ (.CLK(clknet_leaf_63_clk),
    .D(_1244_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ));
 sky130_fd_sc_hd__dfrtp_4 _8250_ (.CLK(clknet_leaf_46_clk),
    .D(_1245_),
    .RESET_B(_0163_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_4 _8251_ (.CLK(clknet_leaf_14_clk),
    .D(_1246_),
    .RESET_B(_0164_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _8252_ (.CLK(clknet_leaf_14_clk),
    .D(_1247_),
    .RESET_B(_0165_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_4 _8253_ (.CLK(clknet_leaf_14_clk),
    .D(_1248_),
    .RESET_B(_0166_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _8254_ (.CLK(clknet_leaf_14_clk),
    .D(_1249_),
    .RESET_B(_0167_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _8255_ (.CLK(clknet_leaf_5_clk),
    .D(_1250_),
    .RESET_B(_0168_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _8256_ (.CLK(clknet_leaf_5_clk),
    .D(_1251_),
    .RESET_B(_0169_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_4 _8257_ (.CLK(clknet_leaf_8_clk),
    .D(_1252_),
    .RESET_B(_0170_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_4 _8258_ (.CLK(clknet_leaf_0_clk),
    .D(_1253_),
    .RESET_B(_0171_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _8259_ (.CLK(clknet_leaf_13_clk),
    .D(_1254_),
    .RESET_B(_0172_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_4 _8260_ (.CLK(clknet_leaf_8_clk),
    .D(_1255_),
    .RESET_B(_0173_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _8261_ (.CLK(clknet_leaf_43_clk),
    .D(_1256_),
    .RESET_B(_0174_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 _8262_ (.CLK(clknet_leaf_10_clk),
    .D(_1257_),
    .RESET_B(_0175_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_4 _8263_ (.CLK(clknet_leaf_13_clk),
    .D(_1258_),
    .RESET_B(_0176_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 _8264_ (.CLK(clknet_leaf_17_clk),
    .D(_1259_),
    .RESET_B(_0177_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _8265_ (.CLK(clknet_leaf_19_clk),
    .D(_1260_),
    .RESET_B(_0178_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _8266_ (.CLK(clknet_leaf_10_clk),
    .D(_1261_),
    .RESET_B(_0179_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_4 _8267_ (.CLK(clknet_leaf_47_clk),
    .D(_1262_),
    .RESET_B(_0180_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _8268_ (.CLK(clknet_leaf_66_clk),
    .D(_1263_),
    .RESET_B(_0181_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_4 _8269_ (.CLK(clknet_leaf_62_clk),
    .D(_1264_),
    .RESET_B(_0182_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_4 _8270_ (.CLK(clknet_leaf_67_clk),
    .D(_1265_),
    .RESET_B(_0183_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_2 _8271_ (.CLK(clknet_leaf_67_clk),
    .D(_1266_),
    .RESET_B(_0184_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 _8272_ (.CLK(clknet_leaf_66_clk),
    .D(_1267_),
    .RESET_B(_0185_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_2 _8273_ (.CLK(clknet_leaf_62_clk),
    .D(_1268_),
    .RESET_B(_0186_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_4 _8274_ (.CLK(clknet_leaf_61_clk),
    .D(_1269_),
    .RESET_B(_0187_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_4 _8275_ (.CLK(clknet_leaf_67_clk),
    .D(_1270_),
    .RESET_B(_0188_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _8276_ (.CLK(clknet_leaf_68_clk),
    .D(_1271_),
    .RESET_B(_0189_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _8277_ (.CLK(clknet_leaf_80_clk),
    .D(_1272_),
    .RESET_B(_0190_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 _8278_ (.CLK(clknet_leaf_79_clk),
    .D(_1273_),
    .RESET_B(_0191_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 _8279_ (.CLK(clknet_leaf_62_clk),
    .D(_1274_),
    .RESET_B(_0192_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_4 _8280_ (.CLK(clknet_leaf_12_clk),
    .D(net707),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8281_ (.CLK(clknet_leaf_12_clk),
    .D(net701),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8282_ (.CLK(clknet_leaf_45_clk),
    .D(net978),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8283_ (.CLK(clknet_leaf_11_clk),
    .D(net1324),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8284_ (.CLK(clknet_leaf_14_clk),
    .D(net2147),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8285_ (.CLK(clknet_leaf_12_clk),
    .D(net2075),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8286_ (.CLK(clknet_leaf_45_clk),
    .D(net577),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8287_ (.CLK(clknet_leaf_4_clk),
    .D(net768),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8288_ (.CLK(clknet_leaf_4_clk),
    .D(net1758),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8289_ (.CLK(clknet_leaf_10_clk),
    .D(net795),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8290_ (.CLK(clknet_leaf_1_clk),
    .D(net1966),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8291_ (.CLK(clknet_leaf_13_clk),
    .D(net2004),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8292_ (.CLK(clknet_leaf_12_clk),
    .D(net627),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8293_ (.CLK(clknet_leaf_43_clk),
    .D(net1811),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8294_ (.CLK(clknet_leaf_10_clk),
    .D(net2014),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8295_ (.CLK(clknet_leaf_13_clk),
    .D(net2013),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8296_ (.CLK(clknet_leaf_17_clk),
    .D(net2072),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8297_ (.CLK(clknet_leaf_44_clk),
    .D(net1034),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8298_ (.CLK(clknet_leaf_10_clk),
    .D(net1948),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8299_ (.CLK(clknet_leaf_47_clk),
    .D(net1973),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8300_ (.CLK(clknet_leaf_66_clk),
    .D(net786),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8301_ (.CLK(clknet_leaf_62_clk),
    .D(net2142),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8302_ (.CLK(clknet_leaf_67_clk),
    .D(net2165),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8303_ (.CLK(clknet_leaf_67_clk),
    .D(net1711),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8304_ (.CLK(clknet_leaf_66_clk),
    .D(net2071),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8305_ (.CLK(clknet_leaf_62_clk),
    .D(net834),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8306_ (.CLK(clknet_leaf_61_clk),
    .D(net2003),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8307_ (.CLK(clknet_leaf_68_clk),
    .D(net2194),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8308_ (.CLK(clknet_leaf_68_clk),
    .D(net2005),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8309_ (.CLK(clknet_leaf_80_clk),
    .D(net1696),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8310_ (.CLK(clknet_leaf_79_clk),
    .D(net2064),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8311_ (.CLK(clknet_leaf_63_clk),
    .D(net2150),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[31] ));
 sky130_fd_sc_hd__ebufn_1 _8319_ (.A(net471),
    .TE_B(_3562_),
    .Z(_0064_));
 sky130_fd_sc_hd__conb_1 _8319__471 (.HI(net471));
 sky130_fd_sc_hd__ebufn_1 _8320_ (.A(net472),
    .TE_B(_3563_),
    .Z(_0065_));
 sky130_fd_sc_hd__conb_1 _8320__472 (.HI(net472));
 sky130_fd_sc_hd__ebufn_1 _8321_ (.A(net466),
    .TE_B(_3564_),
    .Z(_0066_));
 sky130_fd_sc_hd__conb_1 _8321__466 (.LO(net466));
 sky130_fd_sc_hd__ebufn_1 _8322_ (.A(net467),
    .TE_B(_3565_),
    .Z(_0067_));
 sky130_fd_sc_hd__conb_1 _8322__467 (.LO(net467));
 sky130_fd_sc_hd__ebufn_1 _8323_ (.A(net468),
    .TE_B(_3566_),
    .Z(_0068_));
 sky130_fd_sc_hd__conb_1 _8323__468 (.LO(net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__conb_1 core_469 (.LO(net469));
 sky130_fd_sc_hd__conb_1 core_470 (.LO(net470));
 sky130_fd_sc_hd__buf_6 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(_2424_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_6 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(net2046),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net170),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net2046),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 fanout174 (.A(_2423_),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net182),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net182),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_2423_),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_16 fanout184 (.A(_1708_),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(_1435_),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(_1435_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(_1476_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(_1476_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(_1476_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(_1467_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(_1467_),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net201),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_6 fanout201 (.A(_1466_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(net204),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_8 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_1450_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(_1449_),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_8 fanout207 (.A(net209),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(_1434_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net213),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(_1425_),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(_1425_),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net217),
    .X(net215));
 sky130_fd_sc_hd__buf_2 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(_1424_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_8 fanout219 (.A(_2724_),
    .X(net219));
 sky130_fd_sc_hd__buf_6 fanout220 (.A(_2723_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(_2723_),
    .X(net221));
 sky130_fd_sc_hd__buf_8 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_8 fanout223 (.A(_3465_),
    .X(net223));
 sky130_fd_sc_hd__buf_8 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_8 fanout225 (.A(_3461_),
    .X(net225));
 sky130_fd_sc_hd__buf_6 fanout226 (.A(_3457_),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(_3457_),
    .X(net227));
 sky130_fd_sc_hd__buf_6 fanout228 (.A(_3449_),
    .X(net228));
 sky130_fd_sc_hd__buf_6 fanout229 (.A(_3449_),
    .X(net229));
 sky130_fd_sc_hd__buf_6 fanout230 (.A(_3437_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 fanout231 (.A(_3437_),
    .X(net231));
 sky130_fd_sc_hd__buf_8 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_8 fanout233 (.A(_3433_),
    .X(net233));
 sky130_fd_sc_hd__buf_6 fanout234 (.A(_2623_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_8 fanout235 (.A(_2623_),
    .X(net235));
 sky130_fd_sc_hd__buf_6 fanout236 (.A(_2583_),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(_2583_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_16 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_16 fanout239 (.A(_1370_),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout240 (.A(_1368_),
    .X(net240));
 sky130_fd_sc_hd__buf_8 fanout241 (.A(_1368_),
    .X(net241));
 sky130_fd_sc_hd__buf_8 fanout242 (.A(_1352_),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_16 fanout243 (.A(_1352_),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(net248),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(_1324_),
    .X(net248));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_8 fanout250 (.A(_1324_),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(_1324_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_8 fanout254 (.A(net257),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_8 fanout258 (.A(_1323_),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(_1323_),
    .X(net261));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_8 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 fanout264 (.A(_1323_),
    .X(net264));
 sky130_fd_sc_hd__buf_6 fanout265 (.A(_3469_),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_8 fanout266 (.A(_3469_),
    .X(net266));
 sky130_fd_sc_hd__buf_8 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_8 fanout268 (.A(_3463_),
    .X(net268));
 sky130_fd_sc_hd__buf_8 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_8 fanout270 (.A(_3459_),
    .X(net270));
 sky130_fd_sc_hd__buf_8 fanout271 (.A(_3455_),
    .X(net271));
 sky130_fd_sc_hd__buf_8 fanout272 (.A(_3455_),
    .X(net272));
 sky130_fd_sc_hd__buf_6 fanout273 (.A(_3453_),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_8 fanout274 (.A(_3453_),
    .X(net274));
 sky130_fd_sc_hd__buf_6 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_8 fanout276 (.A(_3447_),
    .X(net276));
 sky130_fd_sc_hd__buf_8 fanout277 (.A(_3435_),
    .X(net277));
 sky130_fd_sc_hd__buf_6 fanout278 (.A(_3435_),
    .X(net278));
 sky130_fd_sc_hd__buf_8 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_8 fanout280 (.A(_3431_),
    .X(net280));
 sky130_fd_sc_hd__buf_6 fanout281 (.A(_2719_),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_8 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__buf_6 fanout283 (.A(_2712_),
    .X(net283));
 sky130_fd_sc_hd__buf_8 fanout284 (.A(_2663_),
    .X(net284));
 sky130_fd_sc_hd__buf_8 fanout285 (.A(_2663_),
    .X(net285));
 sky130_fd_sc_hd__buf_8 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_8 fanout287 (.A(_2628_),
    .X(net287));
 sky130_fd_sc_hd__buf_6 fanout288 (.A(_2621_),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_8 fanout289 (.A(_2621_),
    .X(net289));
 sky130_fd_sc_hd__buf_6 fanout290 (.A(_2587_),
    .X(net290));
 sky130_fd_sc_hd__buf_8 fanout291 (.A(_2587_),
    .X(net291));
 sky130_fd_sc_hd__buf_6 fanout292 (.A(_2581_),
    .X(net292));
 sky130_fd_sc_hd__buf_6 fanout293 (.A(_2581_),
    .X(net293));
 sky130_fd_sc_hd__buf_8 fanout294 (.A(_2546_),
    .X(net294));
 sky130_fd_sc_hd__buf_8 fanout295 (.A(_2546_),
    .X(net295));
 sky130_fd_sc_hd__buf_6 fanout296 (.A(_2545_),
    .X(net296));
 sky130_fd_sc_hd__buf_6 fanout297 (.A(_2545_),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_8 fanout298 (.A(_1472_),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_8 fanout299 (.A(_1440_),
    .X(net299));
 sky130_fd_sc_hd__buf_6 fanout300 (.A(_1360_),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 fanout301 (.A(_1360_),
    .X(net301));
 sky130_fd_sc_hd__buf_8 fanout302 (.A(_1344_),
    .X(net302));
 sky130_fd_sc_hd__buf_8 fanout303 (.A(_1335_),
    .X(net303));
 sky130_fd_sc_hd__buf_12 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__buf_12 fanout305 (.A(_1334_),
    .X(net305));
 sky130_fd_sc_hd__buf_6 fanout306 (.A(_3467_),
    .X(net306));
 sky130_fd_sc_hd__buf_6 fanout307 (.A(_3467_),
    .X(net307));
 sky130_fd_sc_hd__buf_6 fanout308 (.A(_3451_),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_8 fanout309 (.A(_3451_),
    .X(net309));
 sky130_fd_sc_hd__buf_6 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_8 fanout311 (.A(_2716_),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(_2714_),
    .X(net312));
 sky130_fd_sc_hd__buf_8 fanout313 (.A(_2709_),
    .X(net313));
 sky130_fd_sc_hd__buf_4 fanout314 (.A(_2709_),
    .X(net314));
 sky130_fd_sc_hd__buf_8 fanout317 (.A(_2661_),
    .X(net317));
 sky130_fd_sc_hd__buf_8 fanout318 (.A(_2661_),
    .X(net318));
 sky130_fd_sc_hd__buf_6 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__buf_8 fanout320 (.A(_2625_),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_8 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_8 fanout322 (.A(_2585_),
    .X(net322));
 sky130_fd_sc_hd__buf_6 fanout323 (.A(_2585_),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 fanout324 (.A(_2585_),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_8 fanout325 (.A(_2579_),
    .X(net325));
 sky130_fd_sc_hd__buf_6 fanout326 (.A(_2579_),
    .X(net326));
 sky130_fd_sc_hd__buf_8 fanout327 (.A(_2511_),
    .X(net327));
 sky130_fd_sc_hd__buf_8 fanout328 (.A(_2511_),
    .X(net328));
 sky130_fd_sc_hd__buf_6 fanout329 (.A(_2510_),
    .X(net329));
 sky130_fd_sc_hd__buf_6 fanout330 (.A(_2510_),
    .X(net330));
 sky130_fd_sc_hd__buf_6 fanout331 (.A(_1356_),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 fanout332 (.A(_1356_),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(_1651_),
    .X(net333));
 sky130_fd_sc_hd__buf_8 fanout334 (.A(_1642_),
    .X(net334));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(_1632_),
    .X(net335));
 sky130_fd_sc_hd__buf_4 fanout336 (.A(_1622_),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(_1613_),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(_1605_),
    .X(net338));
 sky130_fd_sc_hd__buf_4 fanout339 (.A(_1596_),
    .X(net339));
 sky130_fd_sc_hd__buf_4 fanout340 (.A(_1588_),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(_1579_),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(_1569_),
    .X(net342));
 sky130_fd_sc_hd__buf_4 fanout343 (.A(_1561_),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(_1554_),
    .X(net344));
 sky130_fd_sc_hd__buf_4 fanout345 (.A(_1545_),
    .X(net345));
 sky130_fd_sc_hd__buf_4 fanout346 (.A(_1535_),
    .X(net346));
 sky130_fd_sc_hd__buf_4 fanout347 (.A(_1526_),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_8 fanout348 (.A(_1519_),
    .X(net348));
 sky130_fd_sc_hd__buf_4 fanout349 (.A(_1508_),
    .X(net349));
 sky130_fd_sc_hd__buf_4 fanout350 (.A(_1501_),
    .X(net350));
 sky130_fd_sc_hd__buf_4 fanout351 (.A(_1490_),
    .X(net351));
 sky130_fd_sc_hd__buf_4 fanout352 (.A(_1483_),
    .X(net352));
 sky130_fd_sc_hd__buf_4 fanout353 (.A(_1462_),
    .X(net353));
 sky130_fd_sc_hd__buf_4 fanout354 (.A(_1453_),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_8 fanout355 (.A(_1430_),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_8 fanout356 (.A(_1420_),
    .X(net356));
 sky130_fd_sc_hd__buf_4 fanout357 (.A(_1412_),
    .X(net357));
 sky130_fd_sc_hd__buf_4 fanout358 (.A(_1402_),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_8 fanout359 (.A(_1392_),
    .X(net359));
 sky130_fd_sc_hd__buf_4 fanout360 (.A(_1384_),
    .X(net360));
 sky130_fd_sc_hd__buf_4 fanout361 (.A(_1374_),
    .X(net361));
 sky130_fd_sc_hd__buf_8 fanout362 (.A(_1288_),
    .X(net362));
 sky130_fd_sc_hd__buf_6 fanout363 (.A(_1288_),
    .X(net363));
 sky130_fd_sc_hd__buf_12 fanout364 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .X(net364));
 sky130_fd_sc_hd__buf_12 fanout365 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .X(net365));
 sky130_fd_sc_hd__buf_8 fanout366 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .X(net366));
 sky130_fd_sc_hd__buf_8 fanout367 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .X(net367));
 sky130_fd_sc_hd__buf_8 fanout368 (.A(net370),
    .X(net368));
 sky130_fd_sc_hd__buf_8 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_6 fanout370 (.A(net1189),
    .X(net370));
 sky130_fd_sc_hd__buf_8 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_8 fanout372 (.A(net2054),
    .X(net372));
 sky130_fd_sc_hd__buf_8 fanout373 (.A(net375),
    .X(net373));
 sky130_fd_sc_hd__buf_6 fanout374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__buf_4 fanout375 (.A(net2054),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_8 fanout376 (.A(net378),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_4 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_8 fanout378 (.A(net386),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_8 fanout379 (.A(net386),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_4 fanout380 (.A(net386),
    .X(net380));
 sky130_fd_sc_hd__buf_6 fanout381 (.A(net386),
    .X(net381));
 sky130_fd_sc_hd__buf_4 fanout382 (.A(net386),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_8 fanout383 (.A(net386),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_4 fanout384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_8 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_6 fanout386 (.A(net2246),
    .X(net386));
 sky130_fd_sc_hd__buf_8 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_8 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_8 fanout389 (.A(net397),
    .X(net389));
 sky130_fd_sc_hd__buf_8 fanout390 (.A(net397),
    .X(net390));
 sky130_fd_sc_hd__buf_4 fanout391 (.A(net397),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net397),
    .X(net392));
 sky130_fd_sc_hd__buf_4 fanout393 (.A(net397),
    .X(net393));
 sky130_fd_sc_hd__buf_8 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_8 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_8 fanout397 (.A(net1714),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_16 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_8 fanout399 (.A(net2126),
    .X(net399));
 sky130_fd_sc_hd__buf_8 fanout400 (.A(net2233),
    .X(net400));
 sky130_fd_sc_hd__buf_4 fanout401 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net401));
 sky130_fd_sc_hd__buf_8 fanout402 (.A(net2233),
    .X(net402));
 sky130_fd_sc_hd__buf_8 fanout403 (.A(net2233),
    .X(net403));
 sky130_fd_sc_hd__buf_4 fanout404 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_8 fanout405 (.A(net407),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_4 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_8 fanout407 (.A(net415),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_8 fanout408 (.A(net415),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_4 fanout409 (.A(net415),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_8 fanout410 (.A(net415),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(net415),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_8 fanout412 (.A(net415),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_8 fanout414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(net2264),
    .X(net415));
 sky130_fd_sc_hd__buf_8 fanout416 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_4 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_8 fanout418 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net418));
 sky130_fd_sc_hd__buf_8 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_4 fanout420 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net420));
 sky130_fd_sc_hd__buf_8 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_6 fanout422 (.A(net2263),
    .X(net422));
 sky130_fd_sc_hd__buf_6 fanout423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__buf_8 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_8 fanout425 (.A(net2263),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_8 fanout426 (.A(net2095),
    .X(net426));
 sky130_fd_sc_hd__buf_8 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_12 fanout428 (.A(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_4 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_4 fanout430 (.A(net441),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_4 fanout432 (.A(net441),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_8 fanout433 (.A(net441),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_4 fanout434 (.A(net441),
    .X(net434));
 sky130_fd_sc_hd__buf_4 fanout435 (.A(net440),
    .X(net435));
 sky130_fd_sc_hd__buf_4 fanout436 (.A(net440),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_4 fanout437 (.A(net440),
    .X(net437));
 sky130_fd_sc_hd__buf_4 fanout438 (.A(net440),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_4 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_4 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_4 fanout441 (.A(_0069_),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_4 fanout442 (.A(net444),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_8 fanout444 (.A(_0069_),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(_0069_),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(_0069_),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_4 fanout449 (.A(net451),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_8 fanout452 (.A(_0069_),
    .X(net452));
 sky130_fd_sc_hd__buf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_8 fanout454 (.A(net456),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_8 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(_0069_),
    .X(net456));
 sky130_fd_sc_hd__buf_8 fanout457 (.A(net459),
    .X(net457));
 sky130_fd_sc_hd__buf_6 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_4 fanout459 (.A(net63),
    .X(net459));
 sky130_fd_sc_hd__buf_8 fanout460 (.A(net465),
    .X(net460));
 sky130_fd_sc_hd__buf_6 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_4 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(net465),
    .X(net463));
 sky130_fd_sc_hd__buf_6 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_8 fanout465 (.A(net63),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_2 hold1 (.A(net81),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0571_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_0326_),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_0720_),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_0991_),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_0519_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_0350_),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0543_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_0958_),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_1038_),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_1070_),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_1114_),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_1068_),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_0339_),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_0346_),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_1137_),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_1103_),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_0945_),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0547_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_1030_),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_1033_),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_0722_),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_1058_),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_1023_),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_0458_),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_0415_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_0351_),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_0983_),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_0348_),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0525_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_1001_),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_1061_),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_1117_),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_0699_),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_1045_),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_0409_),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_1140_),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_1073_),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_0973_),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_0737_),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0657_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_0334_),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_1150_),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_1108_),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_0292_),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_0256_),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_0969_),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_0955_),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_0623_),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_1076_),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_1097_),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0891_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_1008_),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_0708_),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_0410_),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_0690_),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_0982_),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_1006_),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_1069_),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_0960_),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_1110_),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_0394_),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0669_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_0235_),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_0730_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_1083_),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_0259_),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_0329_),
    .X(net1654));
 sky130_fd_sc_hd__clkbuf_2 hold1119 (.A(net2358),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(_0985_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(_1147_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(_0949_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(_0952_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(_0403_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0536_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(_0428_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(_0244_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(_0255_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(_0702_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(_0407_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(_1080_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(_0943_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(_0391_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(_0453_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(_0408_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0671_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(_0754_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(_0967_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(_0981_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(_0425_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(_1019_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(net119),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_0695_),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_1028_),
    .X(net1700));
 sky130_fd_sc_hd__clkbuf_2 hold1165 (.A(net2360),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(_1116_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(net84),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0563_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_0291_),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_1133_),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_1052_),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(net113),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(_1141_),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(_2436_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_0204_),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_0242_),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_0452_),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_1090_),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_0970_),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0544_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_0941_),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_0290_),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_0477_),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_0364_),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_1127_),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0565_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_1017_),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_0270_),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_0383_),
    .X(net1740));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1205 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(_0947_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(_0254_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0915_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(_0238_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(_1077_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(_0727_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(_0251_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(_0284_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(_0709_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(net128),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_0245_),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_0433_),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_0240_),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0681_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_0249_),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_0283_),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_0261_),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_0447_),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_0281_),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_0424_),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_0260_),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_0713_),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_1016_),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_0371_),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0524_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_0253_),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_0246_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_0439_),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_0443_),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_1078_),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_1000_),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_0267_),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_0446_),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_0950_),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_0266_),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0542_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_0234_),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_0258_),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_0289_),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(net103),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(_0272_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(_0264_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(_0250_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(_0287_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(_0282_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(_0370_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(_0437_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0555_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(_0279_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(_0948_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(_0376_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(_0233_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_0372_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(_0230_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(_0236_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(_0357_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(_0276_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(_0288_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0658_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(_0269_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(_0273_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(_0366_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(_0441_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(_0278_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[25] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(_0445_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(_0412_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(_0386_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(_0431_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(_0252_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_1178_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(_1135_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(_0265_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(_0247_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_0285_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(_0380_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_0237_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(_0435_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_0277_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(_0231_),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(_0436_),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0561_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(_0961_),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(_0426_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_0257_),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(_0434_),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(_0359_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(_0274_),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(_0432_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(_0448_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(_0232_),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(_0280_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0574_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(_0263_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(_0365_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(_0438_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(_0275_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(_0752_),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_0361_),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(_0374_),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(_0268_),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_0442_),
    .X(net1923));
 sky130_fd_sc_hd__clkbuf_4 hold1388 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_2428_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0667_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(_0355_),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(_0381_),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(_0444_),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(_0369_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(_0248_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_1615_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(_0429_),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(_0382_),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(_0377_),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(_0243_),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(_0422_),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0588_),
    .X(net677));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1410 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(_0791_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(net108),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_0286_),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_0379_),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(_0363_),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(_1239_),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_0450_),
    .X(net1958));
 sky130_fd_sc_hd__buf_2 hold1423 (.A(net2357),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(_0449_),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_0430_),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(_0356_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0566_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(net100),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(_0367_),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(_0378_),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_0427_),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(net109),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(_0368_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(_0420_),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(_0384_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(_0373_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(_0423_),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(_0419_),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0537_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(_0360_),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(_0241_),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(_0271_),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(_0385_),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(_0362_),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(_0440_),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(_0375_),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(_0239_),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(net116),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(net101),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(net118),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0678_),
    .X(net683));
 sky130_fd_sc_hd__buf_1 hold1470 (.A(net2364),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ),
    .X(net2007));
 sky130_fd_sc_hd__buf_1 hold1472 (.A(net2361),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(_1527_),
    .X(net2011));
 sky130_fd_sc_hd__buf_1 hold1476 (.A(net2369),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(net105),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(net104),
    .X(net2014));
 sky130_fd_sc_hd__buf_1 hold1479 (.A(net2362),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ),
    .X(net684));
 sky130_fd_sc_hd__buf_1 hold1480 (.A(net2367),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ),
    .X(net2017));
 sky130_fd_sc_hd__buf_4 hold1482 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(_2426_),
    .X(net2019));
 sky130_fd_sc_hd__clkbuf_2 hold1484 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(_2438_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(_0205_),
    .X(net2022));
 sky130_fd_sc_hd__clkbuf_2 hold1487 (.A(net2378),
    .X(net2023));
 sky130_fd_sc_hd__buf_1 hold1488 (.A(net2372),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0675_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_1241_),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ),
    .X(net2027));
 sky130_fd_sc_hd__buf_1 hold1492 (.A(_1927_),
    .X(net2028));
 sky130_fd_sc_hd__buf_2 hold1493 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(_2453_),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(_0213_),
    .X(net2031));
 sky130_fd_sc_hd__buf_2 hold1496 (.A(net2379),
    .X(net2032));
 sky130_fd_sc_hd__buf_1 hold1497 (.A(net2368),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(_0308_),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ),
    .X(net2036));
 sky130_fd_sc_hd__buf_2 hold1501 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ),
    .X(net2037));
 sky130_fd_sc_hd__buf_2 hold1502 (.A(_2037_),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(_0216_),
    .X(net2039));
 sky130_fd_sc_hd__buf_1 hold1504 (.A(net2365),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ),
    .X(net2041));
 sky130_fd_sc_hd__clkbuf_2 hold1506 (.A(net2370),
    .X(net2042));
 sky130_fd_sc_hd__buf_2 hold1507 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_1223_),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\U_CONTROL_UNIT.i_jump_EX ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0554_),
    .X(net687));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1510 (.A(_3471_),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(_0315_),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(_1914_),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ),
    .X(net2053));
 sky130_fd_sc_hd__buf_2 hold1518 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(_2434_),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_4 hold1520 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_2430_),
    .X(net2057));
 sky130_fd_sc_hd__clkbuf_4 hold1522 (.A(net2380),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(_0307_),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(net121),
    .X(net2064));
 sky130_fd_sc_hd__buf_2 hold1529 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0560_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ),
    .X(net2066));
 sky130_fd_sc_hd__buf_1 hold1531 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_1807_),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(_1808_),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_1944_),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(net114),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(net106),
    .X(net2072));
 sky130_fd_sc_hd__buf_1 hold1537 (.A(net2374),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_0314_),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(net125),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_4 hold1540 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .X(net2076));
 sky130_fd_sc_hd__buf_1 hold1541 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(_1743_),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(_1744_),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_1907_),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(_1908_),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ),
    .X(net2082));
 sky130_fd_sc_hd__buf_1 hold1547 (.A(net2371),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(_1394_),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0538_),
    .X(net691));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1550 (.A(net75),
    .X(net2086));
 sky130_fd_sc_hd__clkbuf_2 hold1551 (.A(net2384),
    .X(net2087));
 sky130_fd_sc_hd__buf_1 hold1552 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(_1767_),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_1768_),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(_1921_),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(net70),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(_0262_),
    .X(net2094));
 sky130_fd_sc_hd__buf_2 hold1559 (.A(net2381),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(_0229_),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(_1928_),
    .X(net2099));
 sky130_fd_sc_hd__buf_1 hold1564 (.A(net2376),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_0358_),
    .X(net2102));
 sky130_fd_sc_hd__clkbuf_4 hold1567 (.A(net80),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(_0581_),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0670_),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_2 hold1570 (.A(net2356),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_1815_),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(_1816_),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(_1948_),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_0421_),
    .X(net2112));
 sky130_fd_sc_hd__clkbuf_2 hold1577 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_1728_),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(_1730_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ),
    .X(net694));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1580 (.A(_1897_),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_0583_),
    .X(net2118));
 sky130_fd_sc_hd__clkbuf_2 hold1583 (.A(net2382),
    .X(net2119));
 sky130_fd_sc_hd__buf_1 hold1584 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_1747_),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(_1748_),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(_1909_),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_1911_),
    .X(net2124));
 sky130_fd_sc_hd__clkbuf_2 hold1589 (.A(net2387),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0674_),
    .X(net695));
 sky130_fd_sc_hd__buf_4 hold1590 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(net2126));
 sky130_fd_sc_hd__clkbuf_2 hold1591 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(_2455_),
    .X(net2128));
 sky130_fd_sc_hd__clkbuf_2 hold1593 (.A(net2388),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\U_CONTROL_UNIT.i_branch_EX ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(_1707_),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(net69),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(_1762_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0900_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_1855_),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(_1917_),
    .X(net2137));
 sky130_fd_sc_hd__buf_1 hold1602 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(_1795_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_1796_),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(_1937_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(net111),
    .X(net2142));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1607 (.A(net83),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(_0584_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0682_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(net92),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(net124),
    .X(net2147));
 sky130_fd_sc_hd__buf_2 hold1612 (.A(net2385),
    .X(net2148));
 sky130_fd_sc_hd__clkbuf_2 hold1613 (.A(net2383),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(net122),
    .X(net2150));
 sky130_fd_sc_hd__clkbuf_2 hold1615 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(_1739_),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(_1740_),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(_1905_),
    .X(net2154));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1619 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_1724_),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(_1726_),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(_1894_),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_1719_),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(_1720_),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(_1722_),
    .X(net2162));
 sky130_fd_sc_hd__clkbuf_2 hold1627 (.A(net88),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(net112),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0586_),
    .X(net699));
 sky130_fd_sc_hd__buf_1 hold1630 (.A(net2386),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_1321_),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_1322_),
    .X(net2169));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1634 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net2170));
 sky130_fd_sc_hd__buf_1 hold1635 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(_1926_),
    .X(net2172));
 sky130_fd_sc_hd__buf_1 hold1637 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_1712_),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(_1876_),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_1883_),
    .X(net2176));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1641 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(_1735_),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(_1736_),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_1902_),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ),
    .X(net2181));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1646 (.A(_1598_),
    .X(net2182));
 sky130_fd_sc_hd__buf_1 hold1647 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_1716_),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(_1885_),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_1276_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(net85),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(net68),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(_1799_),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(_1800_),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(_1940_),
    .X(net2191));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1656 (.A(net94),
    .X(net2192));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1657 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(net117),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ),
    .X(net2197));
 sky130_fd_sc_hd__buf_1 hold1662 (.A(net74),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ),
    .X(net2199));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1664 (.A(_1915_),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_1375_),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_1731_),
    .X(net2204));
 sky130_fd_sc_hd__clkbuf_2 hold1669 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0572_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_1782_),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ),
    .X(net2207));
 sky130_fd_sc_hd__buf_2 hold1672 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .X(net2208));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1673 (.A(net184),
    .X(net2209));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1674 (.A(net93),
    .X(net2210));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1675 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(_1786_),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(_1843_),
    .X(net2213));
 sky130_fd_sc_hd__clkbuf_2 hold1678 (.A(_1930_),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_1933_),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(_1715_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(net86),
    .X(net2220));
 sky130_fd_sc_hd__clkbuf_2 hold1685 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ),
    .X(net2221));
 sky130_fd_sc_hd__buf_1 hold1686 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ),
    .X(net2222));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1687 (.A(net71),
    .X(net2223));
 sky130_fd_sc_hd__buf_1 hold1688 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(_1770_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0523_),
    .X(net705));
 sky130_fd_sc_hd__buf_1 hold1690 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(_1880_),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(_1881_),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(_1492_),
    .X(net2232));
 sky130_fd_sc_hd__clkbuf_8 hold1697 (.A(net2327),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(net402),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(_1942_),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ),
    .X(net2239));
 sky130_fd_sc_hd__buf_2 hold1704 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(_1900_),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(_1765_),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(_1919_),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(net120),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_1275_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .X(net2247));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1712 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ),
    .X(net2250));
 sky130_fd_sc_hd__buf_1 hold1715 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .X(net2251));
 sky130_fd_sc_hd__buf_1 hold1716 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(_1699_),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_1702_),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(_2731_),
    .X(net2255));
 sky130_fd_sc_hd__clkbuf_2 hold172 (.A(net2377),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(_0625_),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(_1551_),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(_3159_),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(_0641_),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ),
    .X(net2262));
 sky130_fd_sc_hd__clkbuf_2 hold1727 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0219_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(_1488_),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(_0631_),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(_1923_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ),
    .X(net2272));
 sky130_fd_sc_hd__buf_1 hold1737 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(_1810_),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(_1946_),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ),
    .X(net2279));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1744 (.A(_1643_),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ),
    .X(net2281));
 sky130_fd_sc_hd__buf_1 hold1746 (.A(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(_1819_),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(_1951_),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(_1952_),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0570_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .X(net2290));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1755 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ),
    .X(net2291));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1756 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(_0638_),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(_0642_),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(_1640_),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(_0656_),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .X(net2301));
 sky130_fd_sc_hd__clkbuf_8 hold1766 (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(_1396_),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(_3010_),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0569_),
    .X(net713));
 sky130_fd_sc_hd__buf_1 hold1770 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(_1750_),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(_2910_),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(_1611_),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(_1524_),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0550_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_0640_),
    .X(net2326));
 sky130_fd_sc_hd__buf_1 hold1791 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .X(net2329));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1794 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(_1648_),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(_3309_),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(_0649_),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0535_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(_2819_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(_0627_),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .X(net2343));
 sky130_fd_sc_hd__buf_1 hold1808 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0567_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(net102),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(net110),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(net129),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(net115),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(net127),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(net123),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(net95),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(net67),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(net90),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(net89),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(net126),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0913_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(net79),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(net73),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(net82),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(net91),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(net76),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(net77),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(net78),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(net72),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(net65),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0530_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(net66),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(net87),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(net64),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0622_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0533_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0686_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0562_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0578_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0666_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0573_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0512_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0587_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0580_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0531_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0564_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0922_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0527_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0568_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0549_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0575_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0680_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0904_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0683_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[4] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_1157_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0912_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0553_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0534_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0558_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0579_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net2350),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0867_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0673_),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_2 hold237 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_3439_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0755_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0907_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0684_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0902_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0528_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_0679_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0521_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net2347),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[6] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_1159_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0541_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0881_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0911_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net2348),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0877_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0871_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0924_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_0894_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0910_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0873_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[10] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_1163_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0520_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0914_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0869_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0903_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0893_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0889_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0895_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[5] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_1158_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0866_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0919_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ),
    .X(net565));
 sky130_fd_sc_hd__buf_1 hold290 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_1820_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_1821_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0756_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0906_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0878_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(net2349),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0925_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0883_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0923_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0897_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0870_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0876_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0886_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0908_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0868_),
    .X(net850));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold315 (.A(net2373),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0965_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[29] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_1182_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0668_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0909_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0920_),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 hold324 (.A(net2355),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0917_),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0916_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0872_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_1126_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0885_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_1093_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0896_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0545_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0901_),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0387_),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0892_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0388_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0890_),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0691_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0875_),
    .X(net888));
 sky130_fd_sc_hd__buf_1 hold353 (.A(net2375),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_1231_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0884_),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_1027_),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0879_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0324_),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0887_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[31] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_1184_),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0997_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[3] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_1156_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[13] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_1166_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0693_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0726_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0963_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[28] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_1181_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[16] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0552_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_1169_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_1123_),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_4 hold383 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_8 hold384 (.A(_2036_),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_2435_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0203_),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[23] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_1176_),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_1029_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_1134_),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[27] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_1180_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0723_),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[30] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_1183_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0905_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0661_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0966_),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[17] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_1170_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0964_),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[7] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_1160_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[22] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_1175_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .X(net945));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold41 (.A(net2363),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_1056_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0998_),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_1220_),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_1146_),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[8] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_1161_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[20] ),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_2 hold42 (.A(net2354),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_1173_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0546_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0996_),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0480_),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[9] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_1162_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_8 hold43 (.A(_2425_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_1036_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0732_),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_2 hold433 (.A(net2366),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_0451_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[21] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_1174_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_0888_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0200_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[2] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_1155_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net2245),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0694_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[18] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_1171_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0457_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0481_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_1094_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[12] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_1165_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_0978_),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0719_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0676_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_1092_),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_1057_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0714_),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[14] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_1167_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_1118_),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_1060_),
    .X(net1006));
 sky130_fd_sc_hd__buf_1 hold471 (.A(net2359),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_1012_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0874_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_1107_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0466_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0559_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_1149_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[26] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_1179_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_1054_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_1039_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_1075_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_1087_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0460_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_1138_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_0934_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net107),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0664_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0940_),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0462_),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0418_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0417_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[24] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_1177_),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .X(net1045));
 sky130_fd_sc_hd__buf_2 hold51 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_1132_),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_0933_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0342_),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0389_),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0951_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_2429_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0718_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0454_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0976_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_1053_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0692_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0197_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_1047_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_1105_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_1032_),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0471_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_1085_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_1113_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_1082_),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_1059_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_1049_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[15] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_1168_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0522_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0738_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0402_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0703_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_1031_),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0995_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_1100_),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0465_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_1050_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[11] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_1164_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_1128_),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0529_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_1153_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_1122_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_1120_),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_1041_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0406_),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0744_),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0327_),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_1129_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0469_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_1003_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0685_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0400_),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0739_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_1034_),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0325_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0390_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0880_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0733_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0353_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_1096_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0954_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[19] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_1172_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0659_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0475_),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_1102_),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0456_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_1074_),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0956_),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0323_),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_1111_),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_1043_),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0468_),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0396_),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0548_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0413_),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0340_),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0931_),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_0980_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_1037_),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0987_),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0582_),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_1048_),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0337_),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_0330_),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0532_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_1046_),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_1143_),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_2433_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(_0201_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_1066_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_0345_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(_1104_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(_0977_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(_0751_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(_1099_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_1101_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0540_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_0990_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(_0711_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(_1112_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_0971_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_1055_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_0474_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(_0401_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(_0725_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(_0397_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_0715_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0660_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_0753_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_1010_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_1098_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_1148_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_1018_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(_0942_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_1072_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_0392_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(_1022_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_0946_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0899_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(_0479_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_1004_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(_0743_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_1009_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_1084_),
    .X(net1255));
 sky130_fd_sc_hd__buf_2 hold72 (.A(net2052),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(_1095_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(_0405_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(_0352_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(_0944_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(_1025_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(_0696_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(_0972_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(_0395_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(_0700_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(_1106_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0882_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(_0988_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(_0705_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(_0735_),
    .X(net1281));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold746 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(_0624_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(_1124_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(_0989_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(_0482_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_1065_),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(_0986_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_1044_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0921_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(_0467_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(_0472_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(_0336_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(_0701_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(_0399_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(_0455_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(_0689_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(_1091_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(_0344_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(_0745_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0663_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(_0710_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(_0331_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(_1109_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(_1040_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(net2352),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_0937_),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_0999_),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_0698_),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_0470_),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_0747_),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0672_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0557_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_0354_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_0734_),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_1115_),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_1119_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_0724_),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_0984_),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_1142_),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_0332_),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_0932_),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_0349_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0665_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_0478_),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_0731_),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_0741_),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_1154_),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_0338_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_0729_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_1002_),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_0750_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_0414_),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_0716_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0539_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_0721_),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_1139_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_0939_),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_0968_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_0398_),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_1088_),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_0411_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_0994_),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_1007_),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_1145_),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0577_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_0473_),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_0464_),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_1086_),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_1079_),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_1136_),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_0476_),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_1144_),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_0736_),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_1035_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_0704_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0551_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_0992_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_0740_),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_0938_),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_0979_),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_1125_),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0962_),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_0936_),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_1021_),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_1062_),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_1121_),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0556_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_0343_),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_1005_),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_1081_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_1152_),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_0746_),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net2346),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_1130_),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_1089_),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_1024_),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_0707_),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_0953_),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_1015_),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_1042_),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_0459_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_0461_),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_1014_),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0898_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_0749_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_0393_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_1011_),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_0463_),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_0341_),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_0935_),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_0697_),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_0957_),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_1013_),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_0335_),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0677_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_1026_),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_0328_),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_0975_),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_0717_),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_0333_),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_1131_),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_1063_),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_0416_),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_1020_),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_1151_),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0526_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_0404_),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_0347_),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_0748_),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_0959_),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_0576_),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_0706_),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_0728_),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_0742_),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_0712_),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_0974_),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0662_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_1064_),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_1071_),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_1067_),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_0993_),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_1051_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .X(net1535));
 sky130_fd_sc_hd__buf_1 input1 (.A(i_instr_ID[10]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(i_instr_ID[19]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(i_instr_ID[20]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(i_instr_ID[21]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(i_instr_ID[22]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(i_instr_ID[23]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(i_instr_ID[24]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(i_instr_ID[25]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(i_instr_ID[26]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(i_instr_ID[27]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(i_instr_ID[28]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(i_instr_ID[11]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(i_instr_ID[29]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(i_instr_ID[2]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(i_instr_ID[30]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(i_instr_ID[31]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(i_instr_ID[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(i_instr_ID[4]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_instr_ID[5]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(i_instr_ID[6]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(i_instr_ID[7]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(i_instr_ID[8]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(i_instr_ID[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(i_instr_ID[9]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(i_read_data_M[0]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(i_read_data_M[10]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(i_read_data_M[11]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(i_read_data_M[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(i_read_data_M[13]),
    .X(net35));
 sky130_fd_sc_hd__buf_2 input36 (.A(i_read_data_M[14]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(i_read_data_M[15]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(i_read_data_M[16]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(i_read_data_M[17]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(i_instr_ID[13]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(i_read_data_M[18]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(i_read_data_M[19]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(i_read_data_M[1]),
    .X(net42));
 sky130_fd_sc_hd__buf_4 input43 (.A(i_read_data_M[20]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(i_read_data_M[21]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(i_read_data_M[22]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(i_read_data_M[23]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(i_read_data_M[24]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(i_read_data_M[25]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(i_read_data_M[26]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input5 (.A(i_instr_ID[14]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(i_read_data_M[27]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(i_read_data_M[28]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(i_read_data_M[29]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(i_read_data_M[2]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(i_read_data_M[30]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(i_read_data_M[31]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(i_read_data_M[3]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(i_read_data_M[4]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(i_read_data_M[5]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(i_read_data_M[6]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(i_instr_ID[15]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(i_read_data_M[7]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(i_read_data_M[8]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(i_read_data_M[9]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(rst),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input7 (.A(i_instr_ID[16]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(i_instr_ID[17]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(i_instr_ID[18]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 max_cap190 (.A(_1637_),
    .X(net190));
 sky130_fd_sc_hd__buf_4 max_cap315 (.A(_2708_),
    .X(net315));
 sky130_fd_sc_hd__buf_4 max_cap316 (.A(_2708_),
    .X(net316));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(o_pc_IF[10]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(o_pc_IF[11]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(o_pc_IF[12]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(o_pc_IF[13]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(o_pc_IF[14]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(o_pc_IF[15]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(o_pc_IF[16]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(o_pc_IF[17]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(o_pc_IF[18]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(o_pc_IF[19]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(o_pc_IF[20]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(o_pc_IF[21]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(o_pc_IF[22]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(o_pc_IF[23]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(o_pc_IF[24]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(o_pc_IF[25]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(o_pc_IF[26]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(o_pc_IF[27]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(o_pc_IF[28]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(o_pc_IF[29]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(o_pc_IF[2]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(o_pc_IF[30]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(o_pc_IF[31]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(o_pc_IF[3]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(o_pc_IF[4]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(o_pc_IF[5]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(o_pc_IF[6]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(o_pc_IF[7]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(o_pc_IF[8]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(o_pc_IF[9]));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(o_write_data_M[0]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(o_write_data_M[10]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(o_write_data_M[11]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(o_write_data_M[12]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(o_write_data_M[13]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(o_write_data_M[14]));
 sky130_fd_sc_hd__buf_12 output136 (.A(net136),
    .X(o_write_data_M[15]));
 sky130_fd_sc_hd__buf_12 output137 (.A(net137),
    .X(o_write_data_M[16]));
 sky130_fd_sc_hd__buf_12 output138 (.A(net138),
    .X(o_write_data_M[17]));
 sky130_fd_sc_hd__buf_12 output139 (.A(net139),
    .X(o_write_data_M[18]));
 sky130_fd_sc_hd__buf_12 output140 (.A(net140),
    .X(o_write_data_M[19]));
 sky130_fd_sc_hd__buf_12 output141 (.A(net141),
    .X(o_write_data_M[1]));
 sky130_fd_sc_hd__buf_12 output142 (.A(net142),
    .X(o_write_data_M[20]));
 sky130_fd_sc_hd__buf_12 output143 (.A(net143),
    .X(o_write_data_M[21]));
 sky130_fd_sc_hd__buf_12 output144 (.A(net144),
    .X(o_write_data_M[22]));
 sky130_fd_sc_hd__buf_12 output145 (.A(net145),
    .X(o_write_data_M[23]));
 sky130_fd_sc_hd__buf_12 output146 (.A(net146),
    .X(o_write_data_M[24]));
 sky130_fd_sc_hd__buf_12 output147 (.A(net147),
    .X(o_write_data_M[25]));
 sky130_fd_sc_hd__buf_12 output148 (.A(net148),
    .X(o_write_data_M[26]));
 sky130_fd_sc_hd__buf_12 output149 (.A(net149),
    .X(o_write_data_M[27]));
 sky130_fd_sc_hd__buf_12 output150 (.A(net150),
    .X(o_write_data_M[28]));
 sky130_fd_sc_hd__buf_12 output151 (.A(net151),
    .X(o_write_data_M[29]));
 sky130_fd_sc_hd__buf_12 output152 (.A(net152),
    .X(o_write_data_M[2]));
 sky130_fd_sc_hd__buf_12 output153 (.A(net153),
    .X(o_write_data_M[30]));
 sky130_fd_sc_hd__buf_12 output154 (.A(net154),
    .X(o_write_data_M[31]));
 sky130_fd_sc_hd__buf_12 output155 (.A(net155),
    .X(o_write_data_M[3]));
 sky130_fd_sc_hd__buf_12 output156 (.A(net156),
    .X(o_write_data_M[4]));
 sky130_fd_sc_hd__buf_12 output157 (.A(net157),
    .X(o_write_data_M[5]));
 sky130_fd_sc_hd__buf_12 output158 (.A(net158),
    .X(o_write_data_M[6]));
 sky130_fd_sc_hd__buf_12 output159 (.A(net159),
    .X(o_write_data_M[7]));
 sky130_fd_sc_hd__buf_12 output160 (.A(net160),
    .X(o_write_data_M[8]));
 sky130_fd_sc_hd__buf_12 output161 (.A(net161),
    .X(o_write_data_M[9]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(o_data_addr_M[0]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(o_data_addr_M[10]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(o_data_addr_M[11]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(o_data_addr_M[12]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(o_data_addr_M[13]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(o_data_addr_M[14]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(o_data_addr_M[15]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(o_data_addr_M[16]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(o_data_addr_M[17]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(o_data_addr_M[18]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(o_data_addr_M[19]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(o_data_addr_M[1]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(o_data_addr_M[20]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(o_data_addr_M[21]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(o_data_addr_M[22]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(o_data_addr_M[23]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(o_data_addr_M[24]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(o_data_addr_M[25]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(o_data_addr_M[26]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(o_data_addr_M[27]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(o_data_addr_M[28]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(o_data_addr_M[29]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(o_data_addr_M[2]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(o_data_addr_M[30]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(o_data_addr_M[31]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(o_data_addr_M[3]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(o_data_addr_M[4]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(o_data_addr_M[5]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(o_data_addr_M[6]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(o_data_addr_M[7]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(o_data_addr_M[8]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(o_data_addr_M[9]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(o_funct3_MEM[0]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(o_funct3_MEM[1]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(o_funct3_MEM[2]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(o_mem_write_M));
 sky130_fd_sc_hd__clkbuf_1 wire185 (.A(_3186_),
    .X(net185));
 assign o_pc_IF[0] = net469;
 assign o_pc_IF[1] = net470;
endmodule

