* NGSPICE file created from uart_wbs_bridge.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

.subckt uart_wbs_bridge clk i_start_rx i_uart_rx o_uart_tx rst vccd1 vssd1 wb_ack_i
+ wb_adr_o[0] wb_adr_o[10] wb_adr_o[11] wb_adr_o[12] wb_adr_o[13] wb_adr_o[14] wb_adr_o[15]
+ wb_adr_o[1] wb_adr_o[2] wb_adr_o[3] wb_adr_o[4] wb_adr_o[5] wb_adr_o[6] wb_adr_o[7]
+ wb_adr_o[8] wb_adr_o[9] wb_cyc_o wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12]
+ wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19]
+ wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25]
+ wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31]
+ wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9]
+ wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15]
+ wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21]
+ wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28]
+ wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5]
+ wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_stb_o wb_we_o
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0956__A0 hold55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0759__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1270_ _1340_/CLK _1270_/D _1084_/Y vssd1 vssd1 vccd1 vccd1 _1270_/Q sky130_fd_sc_hd__dfrtp_1
X_0985_ _0985_/A _0985_/B vssd1 vssd1 vccd1 vccd1 _0988_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1399_ _1404_/CLK _1399_/D _1213_/Y vssd1 vssd1 vccd1 vccd1 _1399_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout105 _1197_/A vssd1 vssd1 vccd1 vccd1 _1221_/A sky130_fd_sc_hd__buf_4
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0938__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _1260_/Q vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _1300_/Q vssd1 vssd1 vccd1 vccd1 _0853_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _1000_/X vssd1 vssd1 vccd1 vccd1 _1274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0770_ hold152/X _1374_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 _0770_/X sky130_fd_sc_hd__mux2_1
X_1322_ _1340_/CLK _1322_/D _1136_/Y vssd1 vssd1 vccd1 vccd1 _1322_/Q sky130_fd_sc_hd__dfrtp_1
X_1253_ _1331_/CLK _1253_/D _1067_/Y vssd1 vssd1 vccd1 vccd1 _1253_/Q sky130_fd_sc_hd__dfrtp_1
X_1184_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1184_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1417_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0968_ hold26/X _0958_/X _0967_/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__a21o_1
XFILLER_0_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0899_ _0989_/B _0923_/B _0946_/A2 hold4/X vssd1 vssd1 vccd1 vccd1 _1338_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0822_ _0786_/Y _0803_/X _0821_/X _0796_/Y _0821_/A vssd1 vssd1 vccd1 vccd1 _0822_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0753_ _0752_/Y _0687_/C hold305/X _0684_/X vssd1 vssd1 vccd1 vccd1 _0753_/X sky130_fd_sc_hd__a2bb2o_1
X_0684_ _1048_/A _0684_/B vssd1 vssd1 vccd1 vccd1 _0684_/X sky130_fd_sc_hd__or2_1
X_1305_ _1348_/CLK _1305_/D _1119_/Y vssd1 vssd1 vccd1 vccd1 _1305_/Q sky130_fd_sc_hd__dfrtp_1
X_1236_ _1390_/CLK _1236_/D _1050_/Y vssd1 vssd1 vccd1 vccd1 _1236_/Q sky130_fd_sc_hd__dfrtp_2
X_1167_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1167_/Y sky130_fd_sc_hd__inv_2
X_1098_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1098_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1018__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1021_ hold162/X hold119/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1253_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0805_ _1361_/Q _0813_/C _0807_/B _0815_/A vssd1 vssd1 vccd1 vccd1 _0805_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0771__A1 _1373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0667_ hold48/X hold58/X _0662_/Y hold240/X vssd1 vssd1 vccd1 vccd1 _1413_/D sky130_fd_sc_hd__a31o_1
X_0736_ _1394_/Q _1393_/Q _1392_/Q _0693_/A vssd1 vssd1 vccd1 vccd1 _0736_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1219_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1219_/Y sky130_fd_sc_hd__inv_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _1270_/Q hold140/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0992__A1 hold149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0719_ _1048_/A _0719_/B _1401_/Q _1400_/Q vssd1 vssd1 vccd1 vccd1 _0720_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1031__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 _1271_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[18] sky130_fd_sc_hd__buf_12
Xoutput75 _1281_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput42 _1250_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[13] sky130_fd_sc_hd__buf_12
Xoutput53 hold89/A vssd1 vssd1 vccd1 vccd1 wb_adr_o[9] sky130_fd_sc_hd__buf_12
Xoutput86 _1262_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[9] sky130_fd_sc_hd__buf_12
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1026__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0984_ _0679_/A _0959_/C _0850_/X _0836_/X vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout106 input3/X vssd1 vssd1 vccd1 vccd1 _1197_/A sky130_fd_sc_hd__clkbuf_8
X_1398_ _1404_/CLK _1398_/D _1212_/Y vssd1 vssd1 vccd1 vccd1 _1398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0938__B2 _1374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 _0999_/X vssd1 vssd1 vccd1 vccd1 _1275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _1322_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _1244_/Q vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold171 _1299_/Q vssd1 vssd1 vccd1 vccd1 _0860_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1321_ _1348_/CLK _1321_/D _1135_/Y vssd1 vssd1 vccd1 vccd1 _1321_/Q sky130_fd_sc_hd__dfrtp_1
X_1252_ _1386_/CLK hold62/X _1066_/Y vssd1 vssd1 vccd1 vccd1 _1252_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0903__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1183_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1183_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0960__S0 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0967_ _0958_/X hold97/A _0967_/C vssd1 vssd1 vccd1 vccd1 _0967_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0898_ _0906_/A _0902_/B _0864_/D vssd1 vssd1 vccd1 vccd1 _0923_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0821_ _0821_/A _0821_/B vssd1 vssd1 vccd1 vccd1 _0821_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0752_ _0752_/A _0752_/B vssd1 vssd1 vccd1 vccd1 _0752_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0683_ _0726_/A _0682_/B _1048_/A vssd1 vssd1 vccd1 vccd1 _0720_/A sky130_fd_sc_hd__a21oi_1
X_1166_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1166_/Y sky130_fd_sc_hd__inv_2
X_1304_ _1340_/CLK _1304_/D _1118_/Y vssd1 vssd1 vccd1 vccd1 _1304_/Q sky130_fd_sc_hd__dfrtp_1
X_1235_ _1348_/CLK _1235_/D _1049_/Y vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1097_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1034__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1020_ _1254_/Q hold203/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1020_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_11_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1407_/CLK sky130_fd_sc_hd__clkbuf_8
X_0804_ _0799_/Y _0802_/X _0803_/X _0796_/Y _0802_/A vssd1 vssd1 vccd1 vccd1 _1363_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0735_ _0684_/B _0695_/Y _0734_/X _1048_/A _0734_/A vssd1 vssd1 vccd1 vccd1 _0735_/X
+ sky130_fd_sc_hd__a32o_1
X_0666_ _0656_/A hold57/X _0668_/B _0662_/B hold18/X vssd1 vssd1 vccd1 vccd1 _0666_/X
+ sky130_fd_sc_hd__o41a_1
X_1149_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1149_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1218_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1218_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1029__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1003_ _1271_/Q hold136/X _1003_/S vssd1 vssd1 vccd1 vccd1 _1003_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0718_ _0717_/A _0717_/Y _0718_/S vssd1 vssd1 vccd1 vccd1 _0718_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout100_A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0649_ _0668_/B _0657_/B vssd1 vssd1 vccd1 vccd1 _0649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput65 _1272_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[19] sky130_fd_sc_hd__buf_12
Xoutput87 _1420_/X vssd1 vssd1 vccd1 vccd1 wb_stb_o sky130_fd_sc_hd__buf_12
Xoutput43 _1251_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[14] sky130_fd_sc_hd__buf_12
Xoutput54 _1420_/A vssd1 vssd1 vccd1 vccd1 wb_cyc_o sky130_fd_sc_hd__buf_12
Xoutput76 _1282_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold320 _1320_/Q vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0947__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0983_ hold24/X _0958_/X _0982_/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__a21o_1
Xfanout107 _1162_/A vssd1 vssd1 vccd1 vccd1 _1145_/A sky130_fd_sc_hd__buf_6
X_1397_ _1404_/CLK _1397_/D _1211_/Y vssd1 vssd1 vccd1 vccd1 _1397_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0938__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 _0924_/X vssd1 vssd1 vccd1 vccd1 _1322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _1324_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _0921_/Y vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _1373_/Q vssd1 vssd1 vccd1 vccd1 _0864_/B sky130_fd_sc_hd__buf_2
XANTENNA__1037__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 _1343_/Q vssd1 vssd1 vccd1 vccd1 _0876_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1320_ _1331_/CLK _1320_/D _1134_/Y vssd1 vssd1 vccd1 vccd1 _1320_/Q sky130_fd_sc_hd__dfrtp_1
X_1251_ _1340_/CLK _1251_/D _1065_/Y vssd1 vssd1 vccd1 vccd1 _1251_/Q sky130_fd_sc_hd__dfrtp_1
X_1182_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1182_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0960__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0966_ input32/X input9/X input18/X input26/X _0902_/B _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0967_/C sky130_fd_sc_hd__mux4_1
X_0897_ _0989_/B _0921_/B _0946_/A2 hold180/X vssd1 vssd1 vccd1 vccd1 _1339_/D sky130_fd_sc_hd__a2bb2o_1
X_0820_ _0813_/A _0819_/X _0814_/B vssd1 vssd1 vccd1 vccd1 _0820_/X sky130_fd_sc_hd__o21ba_1
X_0751_ _0745_/A _0749_/X _0750_/X _0749_/B vssd1 vssd1 vccd1 vccd1 _0752_/B sky130_fd_sc_hd__a22o_1
X_1303_ _1340_/CLK _1303_/D _1117_/Y vssd1 vssd1 vccd1 vccd1 _1303_/Q sky130_fd_sc_hd__dfrtp_1
X_0682_ _0726_/A _0682_/B vssd1 vssd1 vccd1 vccd1 _0684_/B sky130_fd_sc_hd__and2_1
X_1165_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1165_/Y sky130_fd_sc_hd__inv_2
X_1096_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1096_/Y sky130_fd_sc_hd__inv_2
X_1234_ _1390_/CLK _1234_/D _0628_/Y vssd1 vssd1 vccd1 vccd1 _1234_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0949_ hold94/X _0957_/S _0931_/Y _0933_/B vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__a22o_1
XANTENNA__0902__B _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0803_ _0823_/D _0803_/B vssd1 vssd1 vccd1 vccd1 _0803_/X sky130_fd_sc_hd__and2_1
X_0665_ hold48/X _0651_/Y _0662_/Y _0664_/X vssd1 vssd1 vccd1 vccd1 _0665_/X sky130_fd_sc_hd__a31o_1
X_0734_ _0734_/A _0734_/B vssd1 vssd1 vccd1 vccd1 _0734_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1079_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1079_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1217_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1217_/Y sky130_fd_sc_hd__inv_2
X_1148_ _1197_/A vssd1 vssd1 vccd1 vccd1 _1148_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__clkbuf_4
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ _1272_/Q hold157/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0910__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0648_ _0632_/A _0668_/A hold48/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__o21a_1
X_0717_ _0717_/A _0762_/S vssd1 vssd1 vccd1 vccd1 _0717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0901__B1 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0717__B _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1404_/CLK sky130_fd_sc_hd__clkbuf_8
Xoutput66 _1254_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput55 _1253_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[0] sky130_fd_sc_hd__buf_12
Xoutput77 _1255_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[2] sky130_fd_sc_hd__buf_12
Xoutput44 _1252_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[15] sky130_fd_sc_hd__buf_12
Xoutput88 _1236_/Q vssd1 vssd1 vccd1 vccd1 wb_we_o sky130_fd_sc_hd__buf_12
XFILLER_0_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold310 _1349_/Q vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _1347_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0982_ _0958_/X hold97/A _0982_/C vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__and3b_1
Xfanout108 input3/X vssd1 vssd1 vccd1 vccd1 _1162_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1396_ _1404_/CLK _1396_/D _1210_/Y vssd1 vssd1 vccd1 vccd1 _1396_/Q sky130_fd_sc_hd__dfrtp_1
Xhold140 _1335_/Q vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _1247_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _1253_/Q vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold195 _1360_/Q vssd1 vssd1 vccd1 vccd1 _0789_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _0920_/X vssd1 vssd1 vccd1 vccd1 _1324_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _0914_/X vssd1 vssd1 vccd1 vccd1 _1328_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1181_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1181_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output54_A _1420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1250_ _1339_/CLK _1250_/D _1064_/Y vssd1 vssd1 vccd1 vccd1 _1250_/Q sky130_fd_sc_hd__dfrtp_1
X_0965_ hold6/X _0958_/X _0964_/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__a21o_1
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0896_ _0906_/A _0902_/B hold149/X vssd1 vssd1 vccd1 vccd1 _0921_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1379_ _1417_/CLK _1379_/D _1193_/Y vssd1 vssd1 vccd1 vccd1 _1379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0750_ hold44/X _1382_/Q hold42/X hold40/X _0692_/S _0749_/A vssd1 vssd1 vccd1 vccd1
+ _0750_/X sky130_fd_sc_hd__mux4_1
X_0681_ _0681_/A _0681_/B _0681_/C _0681_/D vssd1 vssd1 vccd1 vccd1 _0682_/B sky130_fd_sc_hd__or4_1
Xfanout90 _1003_/S vssd1 vssd1 vccd1 vccd1 _1019_/S sky130_fd_sc_hd__buf_6
X_1302_ _1348_/CLK hold95/X _1116_/Y vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfrtp_1
X_1233_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1233_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1164_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1164_/Y sky130_fd_sc_hd__inv_2
X_1095_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1095_/Y sky130_fd_sc_hd__inv_2
X_0948_ hold216/X _0948_/A2 _0929_/Y hold134/X vssd1 vssd1 vccd1 vccd1 _1303_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0879_ _0879_/A hold96/X _0883_/B _0879_/D vssd1 vssd1 vccd1 vccd1 _0879_/Y sky130_fd_sc_hd__nand4_1
X_0802_ _0802_/A _0802_/B vssd1 vssd1 vccd1 vccd1 _0802_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0664_ _0668_/A _0668_/B _0653_/B hold69/X vssd1 vssd1 vccd1 vccd1 _0664_/X sky130_fd_sc_hd__o31a_1
X_0733_ _0733_/A _0733_/B _0733_/C vssd1 vssd1 vccd1 vccd1 _0733_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1216_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1216_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0990__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1147_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1147_/Y sky130_fd_sc_hd__inv_2
X_1078_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1078_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0995__A1 _0864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__buf_2
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0910__B2 _1377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1001_ _1273_/Q hold4/X _1019_/S vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__mux2_1
X_0647_ _0647_/A _0652_/A vssd1 vssd1 vccd1 vccd1 _0657_/B sky130_fd_sc_hd__xor2_1
X_0716_ _0721_/S _0723_/B vssd1 vssd1 vccd1 vccd1 _0718_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0901__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 _1238_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[1] sky130_fd_sc_hd__buf_12
Xoutput67 _1273_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput56 _1263_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xoutput78 _1283_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[30] sky130_fd_sc_hd__buf_12
XANTENNA__0908__B _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold322 _1389_/Q vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold311 _1382_/Q vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 _1390_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0981__S0 hold91/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0972__S0 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0981_ input5/X input35/X input12/X input21/X hold91/A _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0982_/C sky130_fd_sc_hd__mux4_1
XFILLER_0_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout109 input3/X vssd1 vssd1 vccd1 vccd1 _1139_/A sky130_fd_sc_hd__buf_8
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1395_ _1407_/CLK _1395_/D _1209_/Y vssd1 vssd1 vccd1 vccd1 _1395_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0963__S0 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold141 _1004_/X vssd1 vssd1 vccd1 vccd1 _1270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _1304_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _1374_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__buf_1
Xhold152 _1415_/Q vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _1375_/Q vssd1 vssd1 vccd1 vccd1 _0864_/D sky130_fd_sc_hd__clkbuf_2
Xhold185 _1346_/Q vssd1 vssd1 vccd1 vccd1 _0852_/B sky130_fd_sc_hd__buf_2
Xhold196 _0810_/X vssd1 vssd1 vccd1 vccd1 _1360_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0739__A _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1180_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1180_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0964_ _0958_/X hold97/A _0964_/C vssd1 vssd1 vccd1 vccd1 _0964_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_6_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0895_ _0989_/B _0919_/B _0956_/S hold159/X vssd1 vssd1 vccd1 vccd1 _1340_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__0993__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1378_ _1419_/CLK hold68/X _1192_/Y vssd1 vssd1 vccd1 vccd1 _1378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout91 _0948_/A2 vssd1 vssd1 vccd1 vccd1 _0956_/S sky130_fd_sc_hd__buf_4
XFILLER_0_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0680_ _0679_/A _0835_/B _0726_/A vssd1 vssd1 vccd1 vccd1 _1048_/A sky130_fd_sc_hd__a21oi_4
X_1232_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1232_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1301_ _1338_/CLK _1301_/D _1115_/Y vssd1 vssd1 vccd1 vccd1 _1301_/Q sky130_fd_sc_hd__dfrtp_1
X_1094_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1094_/Y sky130_fd_sc_hd__inv_2
X_1163_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1163_/Y sky130_fd_sc_hd__inv_2
XANTENNA_hold91_A hold91/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0947_ hold130/X _0948_/A2 _0927_/Y _0933_/B vssd1 vssd1 vccd1 vccd1 _0947_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0878_ hold96/X _0883_/B _0879_/D _0879_/A vssd1 vssd1 vccd1 vccd1 _0878_/X sky130_fd_sc_hd__a31o_1
XANTENNA__0896__C_N hold149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ _0823_/D _0792_/Y _0800_/X _0796_/Y _0784_/A vssd1 vssd1 vccd1 vccd1 _0801_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0663_ hold48/X _0629_/Y _0662_/Y _0661_/X vssd1 vssd1 vccd1 vccd1 _1415_/D sky130_fd_sc_hd__a31o_1
X_0732_ _0734_/A _1390_/Q _0734_/B _0696_/A vssd1 vssd1 vccd1 vccd1 _0732_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1215_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1215_/Y sky130_fd_sc_hd__inv_2
X_1146_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1146_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1077_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1077_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0910__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1000_ _1274_/Q hold180/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0715_ _0715_/A _1400_/Q _0724_/B vssd1 vssd1 vccd1 vccd1 _0723_/B sky130_fd_sc_hd__and3_1
X_0646_ _0647_/A _0652_/A vssd1 vssd1 vccd1 vccd1 _0662_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1129_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1129_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput46 _1239_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[2] sky130_fd_sc_hd__buf_12
Xoutput57 hold81/A vssd1 vssd1 vccd1 vccd1 wb_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput79 _1284_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xoutput68 _1274_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[21] sky130_fd_sc_hd__buf_12
XFILLER_0_1_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold301 _1357_/Q vssd1 vssd1 vccd1 vccd1 _0814_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _1368_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold323 _1285_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0996__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0629_ _0652_/A hold57/X vssd1 vssd1 vccd1 vccd1 _0629_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0981__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0972__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0980_ hold22/X _0958_/X _0979_/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__a21o_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1394_ _1407_/CLK _1394_/D _1208_/Y vssd1 vssd1 vccd1 vccd1 _1394_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0963__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 _1243_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _1251_/Q vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _0947_/X vssd1 vssd1 vccd1 vccd1 _1304_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _0932_/X vssd1 vssd1 vccd1 vccd1 _1318_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _1297_/Q vssd1 vssd1 vccd1 vccd1 _0859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _0770_/X vssd1 vssd1 vccd1 vccd1 _1374_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _1345_/Q vssd1 vssd1 vccd1 vccd1 _0906_/A sky130_fd_sc_hd__buf_2
Xhold186 _0892_/B vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0894_ _0906_/A hold91/X _0863_/B vssd1 vssd1 vccd1 vccd1 _0919_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0963_ input33/X input10/X input19/X input28/X _0902_/B _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0964_/C sky130_fd_sc_hd__mux4_1
XANTENNA__0831__C _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1377_ _1417_/CLK hold31/X _1191_/Y vssd1 vssd1 vccd1 vccd1 _1377_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout92 _0946_/A2 vssd1 vssd1 vccd1 vccd1 _0948_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1162_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1162_/Y sky130_fd_sc_hd__inv_2
X_1231_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0940__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1300_ _1338_/CLK _1300_/D _1114_/Y vssd1 vssd1 vccd1 vccd1 _1300_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1093_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1093_/Y sky130_fd_sc_hd__inv_2
X_0946_ hold102/X _0946_/A2 _0925_/Y _0933_/B vssd1 vssd1 vccd1 vccd1 _0946_/X sky130_fd_sc_hd__a22o_1
X_0877_ hold96/X _0883_/B _0879_/D vssd1 vssd1 vccd1 vccd1 _0882_/B sky130_fd_sc_hd__nand3_1
XANTENNA_fanout109_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0800_ _1363_/Q _0802_/B _0784_/A vssd1 vssd1 vccd1 vccd1 _0800_/X sky130_fd_sc_hd__a21o_1
X_0731_ _0730_/A _0684_/X _0729_/Y _0730_/Y vssd1 vssd1 vccd1 vccd1 _0731_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0662_ _0668_/B _0662_/B vssd1 vssd1 vccd1 vccd1 _0662_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0913__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1145_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1145_/Y sky130_fd_sc_hd__inv_2
X_1214_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1214_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1076_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1076_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0999__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0929_ _0931_/A _0929_/B vssd1 vssd1 vccd1 vccd1 _0929_/Y sky130_fd_sc_hd__nor2_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__buf_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0645_ _0652_/A _0651_/B vssd1 vssd1 vccd1 vccd1 _0645_/Y sky130_fd_sc_hd__nor2_1
X_0714_ _0726_/A _0734_/B _0714_/C _0714_/D vssd1 vssd1 vccd1 vccd1 _0724_/B sky130_fd_sc_hd__and4_1
X_1059_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1059_/Y sky130_fd_sc_hd__inv_2
X_1128_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1128_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput69 _1275_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput58 _1265_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput47 _1240_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[3] sky130_fd_sc_hd__buf_12
XANTENNA_fanout89_A _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold313 _1367_/Q vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _1372_/Q vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold302 _1408_/Q vssd1 vssd1 vccd1 vccd1 _0692_/S sky130_fd_sc_hd__buf_1
X_0628_ _1231_/A vssd1 vssd1 vccd1 vccd1 _0628_/Y sky130_fd_sc_hd__inv_2
XANTENNA_hold303_A _1420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1393_ _1407_/CLK _1393_/D _1207_/Y vssd1 vssd1 vccd1 vccd1 _1393_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 _1267_/Q vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _1259_/Q vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _0902_/X vssd1 vssd1 vccd1 vccd1 _0927_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _1331_/Q vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _1239_/Q vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _1265_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _1301_/Q vssd1 vssd1 vccd1 vccd1 _0860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _1268_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _1241_/Q vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0893_ _0989_/B hold92/X _0948_/A2 hold85/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0962_ hold16/X _0958_/X _0961_/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__a21o_1
X_1376_ _1417_/CLK hold37/X _1190_/Y vssd1 vssd1 vccd1 vccd1 _1376_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout93 _0957_/S vssd1 vssd1 vccd1 vccd1 _0946_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1092_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1092_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1161_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1161_/Y sky130_fd_sc_hd__inv_2
X_1230_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1230_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0876_ _0876_/A _0902_/B vssd1 vssd1 vccd1 vccd1 _0879_/D sky130_fd_sc_hd__and2_1
X_0945_ hold75/X _0946_/A2 _0923_/Y _0933_/B vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__a22o_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1359_ _1369_/CLK _1359_/D _1173_/Y vssd1 vssd1 vccd1 vccd1 _1359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0922__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0661_ _0653_/A _0632_/A hold239/X hold152/X vssd1 vssd1 vccd1 vccd1 _0661_/X sky130_fd_sc_hd__o31a_1
X_0730_ _0730_/A _0733_/B vssd1 vssd1 vccd1 vccd1 _0730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1213_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1213_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0913__B2 _1374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1144_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1144_/Y sky130_fd_sc_hd__inv_2
X_1075_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1075_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0928_ hold261/X _0956_/S _0927_/Y _0908_/B vssd1 vssd1 vccd1 vccd1 _1320_/D sky130_fd_sc_hd__a22o_1
X_0859_ _0854_/B _0854_/D _0859_/C _0859_/D vssd1 vssd1 vccd1 vccd1 _0859_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0644_ _0647_/A _0632_/A hold239/X hold67/X vssd1 vssd1 vccd1 vccd1 _0644_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0713_ _0701_/A _1048_/A _0684_/B _0712_/Y vssd1 vssd1 vccd1 vccd1 _0713_/X sky130_fd_sc_hd__a22o_1
X_1058_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1058_/Y sky130_fd_sc_hd__inv_2
X_1127_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1127_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput59 _1266_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput48 _1241_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[4] sky130_fd_sc_hd__buf_12
Xoutput37 _1391_/Q vssd1 vssd1 vccd1 vccd1 o_uart_tx sky130_fd_sc_hd__buf_12
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0975__S0 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold314 _1363_/Q vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0627_ input4/X vssd1 vssd1 vccd1 vccd1 _0837_/B sky130_fd_sc_hd__inv_2
Xhold303 _1420_/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0966__S0 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1392_ _1407_/CLK _1392_/D _1206_/Y vssd1 vssd1 vccd1 vccd1 _1392_/Q sky130_fd_sc_hd__dfrtp_1
Xhold144 _0903_/X vssd1 vssd1 vccd1 vccd1 _1336_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _1237_/Q vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 hold319/X vssd1 vssd1 vccd1 vccd1 _0647_/A sky130_fd_sc_hd__buf_2
Xhold133 _1379_/Q vssd1 vssd1 vccd1 vccd1 _0892_/A sky130_fd_sc_hd__clkbuf_2
Xhold100 _1250_/Q vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _1008_/X vssd1 vssd1 vccd1 vccd1 _1266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _1362_/Q vssd1 vssd1 vccd1 vccd1 _0791_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _1308_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _1309_/Q vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _1407_/Q vssd1 vssd1 vccd1 vccd1 _0707_/S sky130_fd_sc_hd__dlygate4sd3_1
X_0961_ _0958_/X hold97/A _0961_/C vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__and3b_1
X_0892_ _0892_/A _0892_/B vssd1 vssd1 vccd1 vccd1 _0957_/S sky130_fd_sc_hd__nand2_1
X_1375_ _1419_/CLK _1375_/D _1189_/Y vssd1 vssd1 vccd1 vccd1 _1375_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0940__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1160_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1160_/Y sky130_fd_sc_hd__inv_2
X_1091_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1091_/Y sky130_fd_sc_hd__inv_2
X_0944_ hold77/X _0948_/A2 _0921_/Y hold134/X vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0875_ _0884_/B _0883_/B _0875_/C vssd1 vssd1 vccd1 vccd1 _0875_/X sky130_fd_sc_hd__and3b_1
X_1358_ _1369_/CLK _1358_/D _1172_/Y vssd1 vssd1 vccd1 vccd1 _1358_/Q sky130_fd_sc_hd__dfrtp_1
X_1289_ _1383_/CLK hold11/X _1103_/Y vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0922__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0660_ hold48/X _0668_/A _0640_/Y _0645_/Y _0659_/X vssd1 vssd1 vccd1 vccd1 _1416_/D
+ sky130_fd_sc_hd__a41o_1
X_1212_ _1218_/A vssd1 vssd1 vccd1 vccd1 _1212_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0913__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1074_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1074_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1143_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1143_/Y sky130_fd_sc_hd__inv_2
X_0927_ _0931_/A _0927_/B vssd1 vssd1 vccd1 vccd1 _0927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout114_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0789_ _0789_/A _1359_/Q _0821_/B _0811_/C vssd1 vssd1 vccd1 vccd1 _0807_/B sky130_fd_sc_hd__and4_1
X_0858_ _0867_/S _0857_/X _1025_/A vssd1 vssd1 vccd1 vccd1 _1348_/D sky130_fd_sc_hd__a21bo_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__buf_2
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0643_ _0643_/A _0763_/B _0803_/B _0823_/D vssd1 vssd1 vccd1 vccd1 _0668_/B sky130_fd_sc_hd__or4b_4
X_0712_ _0712_/A _0712_/B vssd1 vssd1 vccd1 vccd1 _0712_/Y sky130_fd_sc_hd__nor2_1
X_1126_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1126_/Y sky130_fd_sc_hd__inv_2
X_1057_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1057_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0864__B _0864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput38 _1237_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[0] sky130_fd_sc_hd__buf_12
Xoutput49 _1242_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[5] sky130_fd_sc_hd__buf_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0975__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 _1347_/Q vssd1 vssd1 vccd1 vccd1 _0849_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _1321_/Q vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0966__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0626_ _0876_/A vssd1 vssd1 vccd1 vccd1 _0890_/B sky130_fd_sc_hd__inv_2
X_1109_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1109_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1391_ _1404_/CLK _1391_/D _1205_/Y vssd1 vssd1 vccd1 vccd1 _1391_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_9_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold156 _0943_/X vssd1 vssd1 vccd1 vccd1 _1308_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _1041_/X vssd1 vssd1 vccd1 vccd1 _1237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _1316_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _1377_/Q vssd1 vssd1 vccd1 vccd1 _0863_/B sky130_fd_sc_hd__clkbuf_2
Xhold112 _0653_/X vssd1 vssd1 vccd1 vccd1 _0654_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _0933_/B vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__clkbuf_2
Xhold101 _1028_/X vssd1 vssd1 vccd1 vccd1 _1250_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold178 _1294_/Q vssd1 vssd1 vccd1 vccd1 _0854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _0707_/X vssd1 vssd1 vccd1 vccd1 _1407_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0952__A0 hold149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0960_ input34/X input11/X input20/X input29/X _0902_/B _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0961_/C sky130_fd_sc_hd__mux4_1
XFILLER_0_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0891_ _0891_/A _1345_/Q hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__or3_1
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1374_ _1417_/CLK _1374_/D _1188_/Y vssd1 vssd1 vccd1 vccd1 _1374_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0934__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1090_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1090_/Y sky130_fd_sc_hd__inv_2
X_0943_ hold155/X _0948_/A2 _0919_/Y hold134/X vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__a22o_1
X_0874_ _0874_/A _0889_/B vssd1 vssd1 vccd1 vccd1 _0875_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0916__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1357_ _1369_/CLK _1357_/D _1171_/Y vssd1 vssd1 vccd1 vccd1 _1357_/Q sky130_fd_sc_hd__dfrtp_1
X_1288_ _1383_/CLK hold99/X _1102_/Y vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__0883__A _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0907__B1 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1142_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1142_/Y sky130_fd_sc_hd__inv_2
X_1211_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1211_/Y sky130_fd_sc_hd__inv_2
X_1073_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1073_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0926_ hold224/X _0948_/A2 _0925_/Y _0908_/B vssd1 vssd1 vccd1 vccd1 _1321_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0857_ _0857_/A _0871_/D _0857_/C vssd1 vssd1 vccd1 vccd1 _0857_/X sky130_fd_sc_hd__or3_1
X_0788_ _0788_/A _0821_/B _0811_/C vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__and3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _1411_/CLK _1409_/D _1223_/Y vssd1 vssd1 vccd1 vccd1 _1409_/Q sky130_fd_sc_hd__dfrtp_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0904__C_N hold55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0711_ _0719_/B _0701_/C _0701_/A vssd1 vssd1 vccd1 vccd1 _0712_/B sky130_fd_sc_hd__a21oi_1
X_0642_ _0642_/A _0642_/B _0642_/C _0642_/D vssd1 vssd1 vccd1 vccd1 _0642_/X sky130_fd_sc_hd__or4_1
XFILLER_0_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0864__C _0864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1125_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1125_/Y sky130_fd_sc_hd__inv_2
X_1056_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1056_/Y sky130_fd_sc_hd__inv_2
Xoutput39 _1247_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[10] sky130_fd_sc_hd__buf_12
X_0909_ hold104/X _0946_/A2 _0908_/X hold65/X vssd1 vssd1 vccd1 vccd1 _0909_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold316 _1371_/Q vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold305 _1391_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_0625_ _0906_/A vssd1 vssd1 vccd1 vccd1 _0879_/A sky130_fd_sc_hd__inv_2
X_1039_ hold154/X hold130/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1239_/D sky130_fd_sc_hd__mux2_1
X_1108_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1108_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _1390_/CLK _1390_/D _1204_/Y vssd1 vssd1 vccd1 vccd1 _1390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold157 _1337_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _0944_/X vssd1 vssd1 vccd1 vccd1 _1307_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _0655_/X vssd1 vssd1 vccd1 vccd1 _1418_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _0935_/X vssd1 vssd1 vccd1 vccd1 _1316_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _1240_/Q vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _1305_/Q vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _1249_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _0957_/X vssd1 vssd1 vccd1 vccd1 _1294_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1420__A _1420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0890_ hold96/X _0890_/B _0908_/B vssd1 vssd1 vccd1 vccd1 _0989_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1373_ _1419_/CLK hold70/X _1187_/Y vssd1 vssd1 vccd1 vccd1 _1373_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0934__B2 hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout96 hold300/X vssd1 vssd1 vccd1 vccd1 _0726_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0942_ hold166/X _0956_/S _0917_/Y hold134/X vssd1 vssd1 vccd1 vccd1 _1309_/D sky130_fd_sc_hd__a22o_1
X_0873_ _0852_/B _0837_/X _0847_/X wire94/X _0872_/X vssd1 vssd1 vccd1 vccd1 _0883_/B
+ sky130_fd_sc_hd__a2111oi_4
XANTENNA__0916__B2 _0864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1356_ _1369_/CLK _1356_/D _1170_/Y vssd1 vssd1 vccd1 vccd1 _1356_/Q sky130_fd_sc_hd__dfrtp_1
X_1287_ _1411_/CLK hold23/X _1101_/Y vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1072_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1072_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1210_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1210_/Y sky130_fd_sc_hd__inv_2
X_1141_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1141_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0787_ _0816_/S _0814_/A _0813_/A _0821_/A vssd1 vssd1 vccd1 vccd1 _0811_/C sky130_fd_sc_hd__and4_1
X_0925_ _0931_/A _0925_/B vssd1 vssd1 vccd1 vccd1 _0925_/Y sky130_fd_sc_hd__nor2_1
X_0856_ _0884_/B _0856_/B _0856_/C vssd1 vssd1 vccd1 vccd1 _0857_/C sky130_fd_sc_hd__and3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ _1411_/CLK _1408_/D _1222_/Y vssd1 vssd1 vccd1 vccd1 _1408_/Q sky130_fd_sc_hd__dfrtp_2
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1339_ _1339_/CLK _1339_/D _1153_/Y vssd1 vssd1 vccd1 vccd1 _1339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0641_ _0643_/A _0763_/B _0764_/A _0823_/D vssd1 vssd1 vccd1 vccd1 _0657_/A sky130_fd_sc_hd__or4bb_1
X_0710_ _0710_/A _0710_/B vssd1 vssd1 vccd1 vccd1 _0710_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0978__S0 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1124_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1124_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0864__D _0864_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1055_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1055_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0969__S0 hold91/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0908_ _0884_/A _0908_/B vssd1 vssd1 vccd1 vccd1 _0908_/X sky130_fd_sc_hd__and2b_4
X_0839_ hold308/X _0902_/B vssd1 vssd1 vccd1 vccd1 _0989_/A sky130_fd_sc_hd__nand2b_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0624_ _0852_/B vssd1 vssd1 vccd1 vccd1 _0624_/Y sky130_fd_sc_hd__inv_2
Xhold306 _0753_/X vssd1 vssd1 vccd1 vccd1 _1391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _1378_/Q vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1038_ hold168/X hold102/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1240_/D sky130_fd_sc_hd__mux2_1
X_1107_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1107_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 _1002_/X vssd1 vssd1 vccd1 vccd1 _1272_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _1336_/Q vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _1325_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold316/X vssd1 vssd1 vccd1 vccd1 _0864_/C sky130_fd_sc_hd__buf_2
Xhold125 _1029_/X vssd1 vssd1 vccd1 vccd1 _1249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _0946_/X vssd1 vssd1 vccd1 vccd1 _1305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _1261_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1002__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0943__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1148__A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1372_ _1417_/CLK hold19/X _1186_/Y vssd1 vssd1 vccd1 vccd1 _1372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0934__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout97 hold241/X vssd1 vssd1 vccd1 vccd1 _0823_/D sky130_fd_sc_hd__buf_4
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0941_ hold32/X _0948_/A2 _0985_/B _0864_/C vssd1 vssd1 vccd1 vccd1 _1310_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0872_ _0892_/A _0850_/X _0835_/Y _0874_/A vssd1 vssd1 vccd1 vccd1 _0872_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1355_ _1369_/CLK _1355_/D _1169_/Y vssd1 vssd1 vccd1 vccd1 _1355_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0916__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1286_ _1390_/CLK hold25/X _1100_/Y vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfrtp_1
X_1071_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1071_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1140_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1140_/Y sky130_fd_sc_hd__inv_2
X_0924_ hold193/X _0948_/A2 _0923_/Y _0908_/B vssd1 vssd1 vccd1 vccd1 _0924_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0786_ _0821_/A _0821_/B vssd1 vssd1 vccd1 vccd1 _0786_/Y sky130_fd_sc_hd__nand2_1
X_0855_ _0856_/B _0856_/C vssd1 vssd1 vccd1 vccd1 _0985_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ _1338_/CLK _1338_/D _1152_/Y vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfrtp_1
X_1407_ _1407_/CLK _1407_/D _1221_/Y vssd1 vssd1 vccd1 vccd1 _1407_/Q sky130_fd_sc_hd__dfrtp_1
X_1269_ _1383_/CLK hold13/X _1083_/Y vssd1 vssd1 vccd1 vccd1 _1269_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1010__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0640_ _0763_/B _0640_/B vssd1 vssd1 vccd1 vccd1 _0640_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0978__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1054_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1054_/Y sky130_fd_sc_hd__inv_2
X_1123_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1123_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0907_ _0989_/B _0931_/B _0946_/A2 hold12/X vssd1 vssd1 vccd1 vccd1 _1334_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__0969__S1 _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0769_ hold108/X _1375_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 _0769_/X sky130_fd_sc_hd__mux2_1
X_0838_ _0874_/A _0835_/Y _0836_/X _0837_/X vssd1 vssd1 vccd1 vccd1 _1025_/A sky130_fd_sc_hd__a211oi_4
XANTENNA__1005__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0841__D_N _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0623_ _0788_/A vssd1 vssd1 vccd1 vccd1 _0811_/A sky130_fd_sc_hd__inv_2
XFILLER_0_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold307 _1348_/Q vssd1 vssd1 vccd1 vccd1 _0849_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _1376_/Q vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1106_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1106_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1037_ hold121/X hold75/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1241_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0955__A0 _0864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold115 _1314_/Q vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _1333_/Q vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _1380_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _1003_/X vssd1 vssd1 vccd1 vccd1 _1271_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _1340_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _0918_/X vssd1 vssd1 vccd1 vccd1 _1325_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout92_A _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0937__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1371_ _1417_/CLK hold35/X _1185_/Y vssd1 vssd1 vccd1 vccd1 _1371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1013__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout98 hold241/X vssd1 vssd1 vccd1 vccd1 _0813_/C sky130_fd_sc_hd__buf_2
XANTENNA__0762__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0940_ hold53/X _0946_/A2 _0985_/B _1372_/Q vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__a22o_1
X_0871_ _0871_/A _0889_/B _0892_/B _0871_/D vssd1 vssd1 vccd1 vccd1 wire94/A sky130_fd_sc_hd__nor4_1
XFILLER_0_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1159__A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1354_ _1418_/CLK _1354_/D _1168_/Y vssd1 vssd1 vccd1 vccd1 _1354_/Q sky130_fd_sc_hd__dfrtp_1
X_1285_ _1383_/CLK _1285_/D _1099_/Y vssd1 vssd1 vccd1 vccd1 _1285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1008__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0757__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1070_/Y sky130_fd_sc_hd__inv_2
X_0854_ _0859_/D _0854_/B _0859_/C _0854_/D vssd1 vssd1 vccd1 vccd1 _0856_/C sky130_fd_sc_hd__and4b_1
XFILLER_0_11_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0923_ _0931_/A _0923_/B vssd1 vssd1 vccd1 vccd1 _0923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0785_ _0785_/A _0823_/A _0785_/C _0830_/S vssd1 vssd1 vccd1 vccd1 _0821_/B sky130_fd_sc_hd__and4_2
XANTENNA__0770__A1 _1374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1337_ _1341_/CLK _1337_/D _1151_/Y vssd1 vssd1 vccd1 vccd1 _1337_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ _1339_/CLK _1268_/D _1082_/Y vssd1 vssd1 vccd1 vccd1 _1268_/Q sky130_fd_sc_hd__dfrtp_1
X_1406_ _1407_/CLK _1406_/D _1220_/Y vssd1 vssd1 vccd1 vccd1 _1406_/Q sky130_fd_sc_hd__dfrtp_1
X_1199_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1199_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1122_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1122_/Y sky130_fd_sc_hd__inv_2
X_1053_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1053_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0906_ _0906_/A hold91/X _0864_/C vssd1 vssd1 vccd1 vccd1 _0931_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0837_ _0849_/B _0837_/B _0852_/C vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__and3b_2
X_0768_ hold36/X _1376_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__mux2_1
X_0699_ _0734_/B _0714_/C _0714_/D vssd1 vssd1 vccd1 vccd1 _0719_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout105_A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1021__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap95 _0638_/Y vssd1 vssd1 vccd1 vccd1 _0764_/A sky130_fd_sc_hd__clkbuf_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 _1345_/Q vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0622_ _0635_/A vssd1 vssd1 vccd1 vccd1 _0783_/A sky130_fd_sc_hd__inv_2
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 _1369_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_1105_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1105_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1036_ _1242_/Q hold77/X _1041_/S vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__mux2_1
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1016__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold116 _0937_/X vssd1 vssd1 vccd1 vccd1 _1314_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 _0909_/X vssd1 vssd1 vccd1 vccd1 _1333_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _1326_/Q vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 _0762_/X vssd1 vssd1 vccd1 vccd1 _1380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold318/X vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__clkbuf_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1019_ _1255_/Q hold261/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1019_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0937__B2 _1375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0928__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1370_ _1417_/CLK hold80/X _1184_/Y vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout99 hold91/X vssd1 vssd1 vccd1 vccd1 _0902_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0870_ _0884_/B _0867_/S _0869_/X _0868_/Y vssd1 vssd1 vccd1 vccd1 _1346_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1353_ _1418_/CLK _1353_/D _1167_/Y vssd1 vssd1 vccd1 vccd1 _1353_/Q sky130_fd_sc_hd__dfrtp_1
X_1284_ _1419_/CLK _1284_/D _1098_/Y vssd1 vssd1 vccd1 vccd1 _1284_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ _1275_/Q hold159/X _1021_/S vssd1 vssd1 vccd1 vccd1 _0999_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0922_ hold46/X _0948_/A2 hold150/X _0908_/B vssd1 vssd1 vccd1 vccd1 _1323_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0853_ _0860_/D _0853_/B _0860_/C _0853_/D vssd1 vssd1 vccd1 vccd1 _0856_/B sky130_fd_sc_hd__and4b_1
X_0784_ _0784_/A _0802_/A vssd1 vssd1 vccd1 vccd1 _0794_/C sky130_fd_sc_hd__and2_1
X_1405_ _1407_/CLK _1405_/D _1219_/Y vssd1 vssd1 vccd1 vccd1 _1405_/Q sky130_fd_sc_hd__dfrtp_1
Xinput1 i_start_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
X_1336_ _1341_/CLK _1336_/D _1150_/Y vssd1 vssd1 vccd1 vccd1 _1336_/Q sky130_fd_sc_hd__dfrtp_1
X_1267_ _1386_/CLK _1267_/D _1081_/Y vssd1 vssd1 vccd1 vccd1 _1267_/Q sky130_fd_sc_hd__dfrtp_1
X_1198_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1198_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1019__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1121_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1121_/Y sky130_fd_sc_hd__inv_2
X_1052_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1052_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0905_ _0989_/B _0929_/B _0948_/A2 hold140/X vssd1 vssd1 vccd1 vccd1 _1335_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0767_ hold30/X _1377_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__mux2_1
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0836_ _0835_/Y _0836_/B _0874_/A vssd1 vssd1 vccd1 vccd1 _0836_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0698_ _0698_/A _0730_/A vssd1 vssd1 vccd1 vccd1 _0714_/D sky130_fd_sc_hd__and2_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _1340_/CLK _1319_/D _1133_/Y vssd1 vssd1 vccd1 vccd1 _1319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0621_ hold57/X vssd1 vssd1 vccd1 vccd1 _0651_/B sky130_fd_sc_hd__inv_2
Xhold309 _1346_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1035_ hold175/X hold155/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1243_/D sky130_fd_sc_hd__mux2_1
X_1104_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1104_/Y sky130_fd_sc_hd__inv_2
X_0819_ _1355_/Q _0813_/C _0821_/B _0815_/A vssd1 vssd1 vccd1 vccd1 _0819_/X sky130_fd_sc_hd__a31o_1
XANTENNA__1032__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold117 _1312_/Q vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0946__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold128 _1330_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _0916_/X vssd1 vssd1 vccd1 vccd1 _1326_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold106 _1383_/Q vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ _1256_/Q hold224/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1018_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1027__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 _1019_/S vssd1 vssd1 vccd1 vccd1 _1021_/S sky130_fd_sc_hd__buf_6
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1352_ _1418_/CLK _1352_/D _1166_/Y vssd1 vssd1 vccd1 vccd1 _1352_/Q sky130_fd_sc_hd__dfrtp_1
X_1283_ _1338_/CLK _1283_/D _1097_/Y vssd1 vssd1 vccd1 vccd1 _1283_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0998_ _1276_/Q hold85/X _1021_/S vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
XANTENNA__1040__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0921_ _0931_/A _0921_/B vssd1 vssd1 vccd1 vccd1 _0921_/Y sky130_fd_sc_hd__nor2_1
X_0783_ _0783_/A _0815_/A vssd1 vssd1 vccd1 vccd1 _0783_/Y sky130_fd_sc_hd__nor2_1
X_0852_ _0850_/B _0852_/B _0852_/C vssd1 vssd1 vccd1 vccd1 _0871_/D sky130_fd_sc_hd__and3b_1
X_1335_ _1340_/CLK _1335_/D _1149_/Y vssd1 vssd1 vccd1 vccd1 _1335_/Q sky130_fd_sc_hd__dfrtp_1
X_1404_ _1404_/CLK _1404_/D _1218_/Y vssd1 vssd1 vccd1 vccd1 _1404_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1266_ _1340_/CLK _1266_/D _1080_/Y vssd1 vssd1 vccd1 vccd1 _1266_/Q sky130_fd_sc_hd__dfrtp_1
Xinput2 i_uart_rx vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_1197_ _1197_/A vssd1 vssd1 vccd1 vccd1 _1197_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1035__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1051_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1051_/Y sky130_fd_sc_hd__inv_2
X_1120_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1120_/Y sky130_fd_sc_hd__inv_2
X_0904_ _0906_/A hold91/X hold55/X vssd1 vssd1 vccd1 vccd1 _0929_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0766_ hold67/X hold65/X _0773_/S vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0697_ _0734_/B _0714_/C vssd1 vssd1 vccd1 vccd1 _0729_/B sky130_fd_sc_hd__and2_1
X_0835_ _0679_/A _0835_/B vssd1 vssd1 vccd1 vccd1 _0835_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1318_ _1331_/CLK _1318_/D _1132_/Y vssd1 vssd1 vccd1 vccd1 _1318_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _1331_/CLK _1249_/D _1063_/Y vssd1 vssd1 vccd1 vccd1 _1249_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0723__A _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0620_ _0652_/A vssd1 vssd1 vccd1 vccd1 _0656_/A sky130_fd_sc_hd__inv_2
XFILLER_0_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1034_ hold182/X hold166/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1244_/D sky130_fd_sc_hd__mux2_1
X_1103_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1103_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout110_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0818_ _0815_/B _0818_/B vssd1 vssd1 vccd1 vccd1 _1357_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0749_ _0749_/A _0749_/B _0749_/C vssd1 vssd1 vccd1 vccd1 _0749_/X sky130_fd_sc_hd__or3_1
XFILLER_0_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0900__B _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 _0939_/X vssd1 vssd1 vccd1 vccd1 _1312_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _0912_/X vssd1 vssd1 vccd1 vccd1 _1330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold107 _0759_/X vssd1 vssd1 vccd1 vccd1 _1383_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1017_ hold205/X hold193/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1257_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1038__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout90_A _1003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1023__A2 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1420_ _1420_/A vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__buf_1
X_1351_ _1418_/CLK _1351_/D _1165_/Y vssd1 vssd1 vccd1 vccd1 _1351_/Q sky130_fd_sc_hd__dfrtp_1
X_1282_ _1339_/CLK _1282_/D _1096_/Y vssd1 vssd1 vccd1 vccd1 _1282_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0997_ hold265/X _0864_/C _1019_/S vssd1 vssd1 vccd1 vccd1 _1277_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 _1405_/Q vssd1 vssd1 vccd1 vccd1 _0706_/A sky130_fd_sc_hd__dlygate4sd3_1
X_0920_ hold183/X _0956_/S _0919_/Y _0908_/B vssd1 vssd1 vccd1 vccd1 _0920_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0782_ _0640_/Y _0776_/X hold57/X vssd1 vssd1 vccd1 vccd1 _1367_/D sky130_fd_sc_hd__mux2_1
X_0851_ _0892_/A _0850_/X _1025_/C _1025_/A vssd1 vssd1 vccd1 vccd1 _0867_/S sky130_fd_sc_hd__o211a_1
X_1265_ _1331_/CLK _1265_/D _1079_/Y vssd1 vssd1 vccd1 vccd1 _1265_/Q sky130_fd_sc_hd__dfrtp_1
X_1403_ _1404_/CLK _1403_/D _1217_/Y vssd1 vssd1 vccd1 vccd1 _1403_/Q sky130_fd_sc_hd__dfrtp_1
X_1334_ _1386_/CLK _1334_/D _1148_/Y vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfrtp_1
Xinput3 rst vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1196_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1196_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1050_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1050_/Y sky130_fd_sc_hd__inv_2
X_0903_ _0989_/B _0927_/B _0948_/A2 hold136/X vssd1 vssd1 vccd1 vccd1 _0903_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1197__A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0834_ _0852_/C _0871_/A vssd1 vssd1 vccd1 vccd1 _0959_/C sky130_fd_sc_hd__nand2_2
X_0765_ _0773_/S vssd1 vssd1 vccd1 vccd1 _1379_/D sky130_fd_sc_hd__inv_2
X_0696_ _0696_/A _0734_/A vssd1 vssd1 vccd1 vccd1 _0714_/C sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1317_ _1339_/CLK hold66/X _1131_/Y vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfrtp_1
X_1248_ _1390_/CLK hold84/X _1062_/Y vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfrtp_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1179_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1102_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1102_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1033_ _1245_/Q hold32/X _1041_/S vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__mux2_1
X_0817_ _0814_/A _0640_/B _0775_/Y _0814_/B vssd1 vssd1 vccd1 vccd1 _0818_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0748_ hold28/X hold8/X _1408_/Q vssd1 vssd1 vccd1 vccd1 _0749_/C sky130_fd_sc_hd__mux2_1
XANTENNA_fanout103_A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0679_ _0679_/A _0835_/B vssd1 vssd1 vccd1 vccd1 _0704_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 _1416_/Q vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 _1318_/Q vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1258_/Q hold46/X _1021_/S vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1350_ _1369_/CLK _1350_/D _1164_/Y vssd1 vssd1 vccd1 vccd1 _1350_/Q sky130_fd_sc_hd__dfrtp_1
X_1281_ _1407_/CLK _1281_/D _1095_/Y vssd1 vssd1 vccd1 vccd1 _1281_/Q sky130_fd_sc_hd__dfrtp_1
X_0996_ hold250/X hold55/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1278_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold228_A _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 _0709_/Y vssd1 vssd1 vccd1 vccd1 _0710_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold280 _1392_/Q vssd1 vssd1 vccd1 vccd1 _0743_/S sky130_fd_sc_hd__dlygate4sd3_1
X_0850_ _0852_/C _0850_/B _0852_/B vssd1 vssd1 vccd1 vccd1 _0850_/X sky130_fd_sc_hd__or3_2
X_0781_ _0632_/A _0640_/Y _0653_/B _0776_/X _0652_/A vssd1 vssd1 vccd1 vccd1 _1368_/D
+ sky130_fd_sc_hd__a32o_1
X_1402_ _1404_/CLK _1402_/D _1216_/Y vssd1 vssd1 vccd1 vccd1 _1402_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput4 wb_ack_i vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
X_1333_ _1339_/CLK _1333_/D _1147_/Y vssd1 vssd1 vccd1 vccd1 _1333_/Q sky130_fd_sc_hd__dfrtp_1
X_1264_ _1338_/CLK hold82/X _1078_/Y vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1195_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1195_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0979_ _0958_/X hold97/A _0979_/C vssd1 vssd1 vccd1 vccd1 _0979_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0902_ _0906_/A _0902_/B _1373_/Q vssd1 vssd1 vccd1 vccd1 _0902_/X sky130_fd_sc_hd__or3b_1
X_0833_ _0852_/B _0850_/B _0852_/C vssd1 vssd1 vccd1 vccd1 _0874_/A sky130_fd_sc_hd__and3b_2
X_0764_ _0764_/A _0764_/B vssd1 vssd1 vccd1 vccd1 _0773_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0695_ _0734_/A _0734_/B vssd1 vssd1 vccd1 vccd1 _0695_/Y sky130_fd_sc_hd__nand2_1
X_1178_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1178_/Y sky130_fd_sc_hd__inv_2
X_1247_ _1341_/CLK _1247_/D _1061_/Y vssd1 vssd1 vccd1 vccd1 _1247_/Q sky130_fd_sc_hd__dfrtp_1
X_1316_ _1340_/CLK _1316_/D _1130_/Y vssd1 vssd1 vccd1 vccd1 _1316_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0991__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1101_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1101_/Y sky130_fd_sc_hd__inv_2
X_1032_ hold89/X hold53/X _1041_/S vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__mux2_1
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0816_ _0815_/B _0815_/Y _0816_/S vssd1 vssd1 vccd1 vccd1 _0816_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0747_ _0749_/B _0747_/B vssd1 vssd1 vccd1 vccd1 _0752_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0678_ _0726_/A _0678_/B _0678_/C vssd1 vssd1 vccd1 vccd1 _0678_/X sky130_fd_sc_hd__and3_1
Xhold109 _0769_/X vssd1 vssd1 vccd1 vccd1 _1375_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1015_ hold198/X hold183/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1259_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ _1340_/CLK _1280_/D _1094_/Y vssd1 vssd1 vccd1 vccd1 _1280_/Q sky130_fd_sc_hd__dfrtp_1
X_0995_ hold259/X _0864_/B _1019_/S vssd1 vssd1 vccd1 vccd1 _1279_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0994__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 _1409_/Q vssd1 vssd1 vccd1 vccd1 _0749_/B sky130_fd_sc_hd__clkbuf_2
Xhold281 _0743_/X vssd1 vssd1 vccd1 vccd1 _1392_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _0710_/Y vssd1 vssd1 vccd1 vccd1 _1405_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0780_ _0647_/A _0779_/Y _0777_/X vssd1 vssd1 vccd1 vccd1 _1369_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ _1404_/CLK _1401_/D _1215_/Y vssd1 vssd1 vccd1 vccd1 _1401_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0912__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1332_ _1386_/CLK hold64/X _1146_/Y vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfrtp_1
X_1263_ _1404_/CLK hold72/X _1077_/Y vssd1 vssd1 vccd1 vccd1 _1263_/Q sky130_fd_sc_hd__dfrtp_1
X_1194_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1194_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0978_ input16/X input36/X input13/X input22/X _0902_/B _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0979_/C sky130_fd_sc_hd__mux4_1
XANTENNA__0903__B1 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0901_ _0989_/B _0925_/B _0948_/A2 hold157/X vssd1 vssd1 vccd1 vccd1 _1337_/D sky130_fd_sc_hd__a2bb2o_1
X_0763_ _0823_/D _0763_/B vssd1 vssd1 vccd1 vccd1 _0764_/B sky130_fd_sc_hd__and2_2
XFILLER_0_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0832_ _0852_/B _0850_/B vssd1 vssd1 vccd1 vccd1 _0871_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1315_ _1339_/CLK hold74/X _1129_/Y vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfrtp_1
X_0694_ _0734_/B vssd1 vssd1 vccd1 vccd1 _0694_/Y sky130_fd_sc_hd__inv_2
X_1177_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1177_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1246_ _1390_/CLK hold90/X _1060_/Y vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1390_/CLK sky130_fd_sc_hd__clkbuf_8
X_1031_ hold151/X hold117/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1247_/D sky130_fd_sc_hd__mux2_1
X_1100_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1100_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0815_ _0815_/A _0815_/B vssd1 vssd1 vccd1 vccd1 _0815_/Y sky130_fd_sc_hd__nor2_1
X_0746_ _0692_/S hold126/X _0745_/Y _0744_/X _0749_/A vssd1 vssd1 vccd1 vccd1 _0747_/B
+ sky130_fd_sc_hd__a32o_1
Xinput30 wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0677_ _0726_/A _0678_/C vssd1 vssd1 vccd1 vccd1 _0687_/C sky130_fd_sc_hd__nand2_1
X_1229_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1229_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1014_ hold170/X hold147/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1260_/D sky130_fd_sc_hd__mux2_1
XANTENNA__0997__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0729_ _1048_/A _0729_/B vssd1 vssd1 vccd1 vccd1 _0729_/Y sky130_fd_sc_hd__nand2b_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0767__A1 _1377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0994_ hold276/X hold163/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1280_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0997__A1 _0864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold260 _1282_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _0691_/X vssd1 vssd1 vccd1 vccd1 _1409_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _1401_/Q vssd1 vssd1 vccd1 vccd1 _0715_/A sky130_fd_sc_hd__buf_1
Xhold293 _1397_/Q vssd1 vssd1 vccd1 vccd1 _0696_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1331_ _1331_/CLK _1331_/D _1145_/Y vssd1 vssd1 vccd1 vccd1 _1331_/Q sky130_fd_sc_hd__dfrtp_1
X_1400_ _1404_/CLK _1400_/D _1214_/Y vssd1 vssd1 vccd1 vccd1 _1400_/Q sky130_fd_sc_hd__dfrtp_1
Xinput6 wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0912__B2 _1375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1193_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1193_/Y sky130_fd_sc_hd__inv_2
X_1262_ _1339_/CLK hold3/X _1076_/Y vssd1 vssd1 vccd1 vccd1 _1262_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0977_ hold20/X _0958_/X hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__a21o_1
XFILLER_0_14_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ _0906_/A _0902_/B hold163/X vssd1 vssd1 vccd1 vccd1 _0925_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_51_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0693_ _0693_/A _0740_/S _0742_/S _0743_/S vssd1 vssd1 vccd1 vccd1 _0734_/B sky130_fd_sc_hd__and4_2
X_0762_ hold126/X hold24/X _0762_/S vssd1 vssd1 vccd1 vccd1 _0762_/X sky130_fd_sc_hd__mux2_1
X_0831_ _0906_/A _0876_/A _0902_/B hold96/X vssd1 vssd1 vccd1 vccd1 _0836_/B sky130_fd_sc_hd__or4b_1
X_1314_ _1331_/CLK _1314_/D _1128_/Y vssd1 vssd1 vccd1 vccd1 _1314_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0897__B1 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1176_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1176_/Y sky130_fd_sc_hd__inv_2
X_1245_ _1418_/CLK hold33/X _1059_/Y vssd1 vssd1 vccd1 vccd1 _1245_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1030_ hold83/X hold51/X _1041_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
X_0814_ _0814_/A _0814_/B vssd1 vssd1 vccd1 vccd1 _0815_/B sky130_fd_sc_hd__and2_1
Xinput31 wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
Xinput20 wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_0676_ _0681_/A _0681_/B _0681_/C _0681_/D vssd1 vssd1 vccd1 vccd1 _0678_/C sky130_fd_sc_hd__nor4_1
X_0745_ _0745_/A _1410_/Q vssd1 vssd1 vccd1 vccd1 _0745_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1228_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1228_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1159_ _1197_/A vssd1 vssd1 vccd1 vccd1 _1159_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ hold169/X hold138/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1261_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0659_ _0653_/A _0652_/A _0651_/B _0657_/A hold108/X vssd1 vssd1 vccd1 vccd1 _0659_/X
+ sky130_fd_sc_hd__o41a_1
X_0728_ _0728_/A _0728_/B vssd1 vssd1 vccd1 vccd1 _0728_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout101_A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1411_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__0898__C_N _0864_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0862__A _1375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0993_ hold251/X _0864_/D _1021_/S vssd1 vssd1 vccd1 vccd1 _1281_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold250 _1278_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold283 _0722_/Y vssd1 vssd1 vccd1 vccd1 _0723_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _0732_/X vssd1 vssd1 vccd1 vccd1 _0733_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hold320/X vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__buf_1
Xhold272 hold323/X vssd1 vssd1 vccd1 vccd1 _0679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1330_ _1331_/CLK _1330_/D _1144_/Y vssd1 vssd1 vccd1 vccd1 _1330_/Q sky130_fd_sc_hd__dfrtp_1
X_1261_ _1411_/CLK _1261_/D _1075_/Y vssd1 vssd1 vccd1 vccd1 _1261_/Q sky130_fd_sc_hd__dfrtp_1
Xinput7 wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
X_1192_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1192_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ _0958_/X hold97/X _0976_/C vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__and3b_1
XFILLER_0_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _0823_/D _0796_/Y _0830_/S vssd1 vssd1 vccd1 vccd1 _1351_/D sky130_fd_sc_hd__mux2_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0761_ hold44/X hold22/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__mux2_1
X_0692_ _0720_/A _0687_/C _0692_/S vssd1 vssd1 vccd1 vccd1 _1408_/D sky130_fd_sc_hd__mux2_1
X_1244_ _1331_/CLK _1244_/D _1058_/Y vssd1 vssd1 vccd1 vccd1 _1244_/Q sky130_fd_sc_hd__dfrtp_1
X_1313_ _1390_/CLK hold52/X _1127_/Y vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfrtp_1
X_1175_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1175_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0959_ _1345_/Q hold96/X _0959_/C vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__nor3_4
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
Xinput21 wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
X_0813_ _0813_/A _0821_/A _0813_/C _0821_/B vssd1 vssd1 vccd1 vccd1 _0814_/B sky130_fd_sc_hd__and4_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput32 wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_1
XFILLER_0_16_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0744_ hold106/X hold87/X _1408_/Q vssd1 vssd1 vccd1 vccd1 _0744_/X sky130_fd_sc_hd__mux2_1
X_0675_ _0696_/A _0693_/A _0740_/S _0734_/A vssd1 vssd1 vccd1 vccd1 _0681_/D sky130_fd_sc_hd__or4bb_1
X_1227_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1227_/Y sky130_fd_sc_hd__inv_2
X_1158_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1158_/Y sky130_fd_sc_hd__inv_2
X_1089_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1089_/Y sky130_fd_sc_hd__inv_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1012_ _1262_/Q hold2/X _1019_/S vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0727_ _0730_/A _0726_/A _0729_/B _0698_/A vssd1 vssd1 vccd1 vccd1 _0727_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0658_ hold48/X hold36/X hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0862__B _1373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0992_ hold260/X hold149/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1282_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_7_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1341_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__0915__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 _0666_/X vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _1281_/Q vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _1019_/X vssd1 vssd1 vccd1 vccd1 _1255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _0723_/Y vssd1 vssd1 vccd1 vccd1 _1401_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _0733_/X vssd1 vssd1 vccd1 vccd1 _1397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _0984_/X vssd1 vssd1 vccd1 vccd1 _1285_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1260_ _1340_/CLK _1260_/D _1074_/Y vssd1 vssd1 vccd1 vccd1 _1260_/Q sky130_fd_sc_hd__dfrtp_1
X_1191_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1191_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0975_ input27/X input6/X input14/X input23/X _0902_/B _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0976_/C sky130_fd_sc_hd__mux4_1
X_1389_ _1419_/CLK hold1/X _1203_/Y vssd1 vssd1 vccd1 vccd1 _1389_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ hold311/X hold20/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0691_ _0687_/C _0690_/Y _0684_/X _0749_/B vssd1 vssd1 vccd1 vccd1 _0691_/X sky130_fd_sc_hd__a2bb2o_1
X_1174_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1174_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1243_ _1340_/CLK _1243_/D _1057_/Y vssd1 vssd1 vccd1 vccd1 _1243_/Q sky130_fd_sc_hd__dfrtp_1
X_1312_ _1341_/CLK _1312_/D _1126_/Y vssd1 vssd1 vccd1 vccd1 _1312_/Q sky130_fd_sc_hd__dfrtp_1
X_0889_ _0892_/A _0889_/B vssd1 vssd1 vccd1 vccd1 _0908_/B sky130_fd_sc_hd__and2_4
XFILLER_0_6_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0958_ _0959_/C _0850_/X _0872_/X vssd1 vssd1 vccd1 vccd1 _0958_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0812_ _0811_/A _0809_/X _0811_/X _0823_/D vssd1 vssd1 vccd1 vccd1 _1359_/D sky130_fd_sc_hd__a2bb2o_1
Xinput11 wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
X_0743_ _0726_/A _1048_/A _0743_/S vssd1 vssd1 vccd1 vccd1 _0743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0674_ _0715_/A _0725_/S _0698_/A _0730_/A vssd1 vssd1 vccd1 vccd1 _0681_/C sky130_fd_sc_hd__or4b_1
X_1226_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1226_/Y sky130_fd_sc_hd__inv_2
X_1157_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1157_/Y sky130_fd_sc_hd__inv_2
X_1088_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1088_/Y sky130_fd_sc_hd__inv_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1011_ _1263_/Q hold71/X _1019_/S vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0726_ _0726_/A _0729_/B vssd1 vssd1 vccd1 vccd1 _0733_/B sky130_fd_sc_hd__nand2_1
X_0657_ _0657_/A _0657_/B hold58/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__or3b_1
X_1209_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1209_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0709_ _0726_/A _0712_/A _0733_/A _0706_/A vssd1 vssd1 vccd1 vccd1 _0709_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0924__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ hold256/X _0863_/B _1019_/S vssd1 vssd1 vccd1 vccd1 _1283_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0915__B2 hold55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold285 _1351_/Q vssd1 vssd1 vccd1 vccd1 _0830_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _1350_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _0665_/X vssd1 vssd1 vccd1 vccd1 _1414_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _1402_/Q vssd1 vssd1 vccd1 vccd1 _0721_/S sky130_fd_sc_hd__buf_1
Xhold263 _1410_/Q vssd1 vssd1 vccd1 vccd1 _0749_/A sky130_fd_sc_hd__clkbuf_2
Xhold274 _1411_/Q vssd1 vssd1 vccd1 vccd1 _0745_/A sky130_fd_sc_hd__buf_1
Xhold296 _1234_/Q vssd1 vssd1 vccd1 vccd1 _0835_/B sky130_fd_sc_hd__buf_2
XFILLER_0_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1190_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1190_/Y sky130_fd_sc_hd__inv_2
Xinput9 wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
X_0974_ hold10/X _0958_/X _0973_/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__a21o_1
X_1388_ _1411_/CLK hold9/X _1202_/Y vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1348_/CLK sky130_fd_sc_hd__clkbuf_8
X_0690_ _0690_/A _0690_/B vssd1 vssd1 vccd1 vccd1 _0690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1311_ _1390_/CLK hold54/X _1125_/Y vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfrtp_1
X_1173_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1173_/Y sky130_fd_sc_hd__inv_2
X_1242_ _1418_/CLK hold78/X _1056_/Y vssd1 vssd1 vccd1 vccd1 _1242_/Q sky130_fd_sc_hd__dfrtp_2
X_0957_ _0864_/C _0854_/D _0957_/S vssd1 vssd1 vccd1 vccd1 _0957_/X sky130_fd_sc_hd__mux2_1
X_0888_ _0883_/X _0888_/B vssd1 vssd1 vccd1 vccd1 _1342_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
X_0811_ _0811_/A _0821_/B _0811_/C vssd1 vssd1 vccd1 vccd1 _0811_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput34 wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput23 wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
X_0673_ _0707_/S _0673_/B _0742_/S _0743_/S vssd1 vssd1 vccd1 vccd1 _0681_/B sky130_fd_sc_hd__or4bb_1
X_0742_ _0741_/X _0739_/Y _0742_/S vssd1 vssd1 vccd1 vccd1 _0742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1225_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1225_/Y sky130_fd_sc_hd__inv_2
X_1087_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1087_/Y sky130_fd_sc_hd__inv_2
X_1156_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1156_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ hold81/X hold38/X _1019_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
X_0656_ _0656_/A hold57/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__nor2_1
X_0725_ _0724_/B _0728_/A _0725_/S vssd1 vssd1 vccd1 vccd1 _0725_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0876__B _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1208_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1208_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1139_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0639_ _0823_/D _0764_/A vssd1 vssd1 vccd1 vccd1 _0640_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0708_ _0673_/B _0710_/A _0705_/Y vssd1 vssd1 vccd1 vccd1 _0708_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0924__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0990_ hold247/X hold65/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1284_/D sky130_fd_sc_hd__mux2_1
XANTENNA__0915__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold231 _1365_/Q vssd1 vssd1 vccd1 vccd1 _0794_/A sky130_fd_sc_hd__buf_1
XFILLER_0_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold242 hold321/X vssd1 vssd1 vccd1 vccd1 _0850_/B sky130_fd_sc_hd__buf_2
Xhold253 _0721_/X vssd1 vssd1 vccd1 vccd1 _1402_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 _0708_/X vssd1 vssd1 vccd1 vccd1 _1406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _0688_/X vssd1 vssd1 vccd1 vccd1 _1410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _1403_/Q vssd1 vssd1 vccd1 vccd1 _0700_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold275 _0686_/X vssd1 vssd1 vccd1 vccd1 _1411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _1045_/X vssd1 vssd1 vccd1 vccd1 _1234_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0973_ _0958_/X hold97/A _0973_/C vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__and3b_1
X_1387_ _1411_/CLK hold29/X _1201_/Y vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1000__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1310_ _1341_/CLK _1310_/D _1124_/Y vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfrtp_1
X_1241_ _1338_/CLK _1241_/D _1055_/Y vssd1 vssd1 vccd1 vccd1 _1241_/Q sky130_fd_sc_hd__dfrtp_2
X_1172_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1172_/Y sky130_fd_sc_hd__inv_2
X_0956_ hold55/X _0859_/C _0956_/S vssd1 vssd1 vccd1 vccd1 _1295_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0887_ _0850_/B _0883_/B _0902_/B vssd1 vssd1 vccd1 vccd1 _0888_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0810_ _0813_/C _0807_/B _0809_/X _0789_/A vssd1 vssd1 vccd1 vccd1 _0810_/X sky130_fd_sc_hd__o2bb2a_1
Xinput13 wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
Xinput35 wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput24 wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
X_0672_ _0706_/A _0700_/A _0721_/S _0701_/A vssd1 vssd1 vccd1 vccd1 _0681_/A sky130_fd_sc_hd__or4bb_1
X_0741_ _1392_/Q _1390_/Q vssd1 vssd1 vccd1 vccd1 _0741_/X sky130_fd_sc_hd__and2_1
XFILLER_0_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1224_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1224_/Y sky130_fd_sc_hd__inv_2
X_1086_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1086_/Y sky130_fd_sc_hd__inv_2
X_1155_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1155_/Y sky130_fd_sc_hd__inv_2
X_0939_ hold117/X _0948_/A2 _0985_/B _1373_/Q vssd1 vssd1 vccd1 vccd1 _0939_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0963__A0 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1340_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA_hold174_A _1375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0655_ hold48/X hold30/X _0655_/S vssd1 vssd1 vccd1 vccd1 _0655_/X sky130_fd_sc_hd__mux2_1
X_0724_ _0762_/S _0724_/B vssd1 vssd1 vccd1 vccd1 _0728_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1207_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1207_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1138_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1138_/Y sky130_fd_sc_hd__inv_2
X_1069_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1069_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0936__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0707_ _0702_/X _0705_/Y _0707_/S vssd1 vssd1 vccd1 vccd1 _0707_/X sky130_fd_sc_hd__mux2_1
X_0638_ _0642_/A _0638_/B _0638_/C _0642_/D vssd1 vssd1 vccd1 vccd1 _0638_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__1003__S _1003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0909__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0906__C_N _0864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold243 _1361_/Q vssd1 vssd1 vccd1 vccd1 _0807_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold210 _1364_/Q vssd1 vssd1 vccd1 vccd1 _0784_/A sky130_fd_sc_hd__buf_1
Xhold232 _0798_/X vssd1 vssd1 vccd1 vccd1 _1365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _1280_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _1238_/Q vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold265 _1277_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _0718_/X vssd1 vssd1 vccd1 vccd1 _1403_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _1396_/Q vssd1 vssd1 vccd1 vccd1 _0734_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold298 _1359_/Q vssd1 vssd1 vccd1 vccd1 _0788_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0972_ input30/X input7/X input15/X input24/X _0902_/B _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0973_/C sky130_fd_sc_hd__mux4_1
XFILLER_0_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1386_ _1386_/CLK hold41/X _1200_/Y vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1171_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1171_/Y sky130_fd_sc_hd__inv_2
X_1240_ _1348_/CLK _1240_/D _1054_/Y vssd1 vssd1 vccd1 vccd1 _1240_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0985__B _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0955_ _0864_/B _0854_/B _0956_/S vssd1 vssd1 vccd1 vccd1 _1296_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0886_ _0883_/B _0885_/X _0883_/X _0876_/A vssd1 vssd1 vccd1 vccd1 _1343_/D sky130_fd_sc_hd__o2bb2a_1
XANTENNA__0990__A1 hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1369_ _1369_/CLK _1369_/D _1183_/Y vssd1 vssd1 vccd1 vccd1 _1369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1011__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XANTENNA__0760__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput14 wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
X_0740_ _0739_/B _0739_/Y _0740_/S vssd1 vssd1 vccd1 vccd1 _0740_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0972__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0671_ _0749_/A _0749_/B _1408_/Q vssd1 vssd1 vccd1 vccd1 _0678_/B sky130_fd_sc_hd__and3_1
X_1154_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1154_/Y sky130_fd_sc_hd__inv_2
X_1223_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1223_/Y sky130_fd_sc_hd__inv_2
X_1085_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1085_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0869_ _0859_/X _0860_/X _0985_/A vssd1 vssd1 vccd1 vccd1 _0869_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__0963__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0938_ hold51/X _0946_/A2 _0985_/B _1374_/Q vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__a22o_1
XFILLER_0_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold167_A _1377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1006__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0755__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0723_ _0762_/S _0723_/B _0723_/C vssd1 vssd1 vccd1 vccd1 _0723_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0654_ _0657_/A _0654_/B vssd1 vssd1 vccd1 vccd1 _0655_/S sky130_fd_sc_hd__or2_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1137_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1137_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_7_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1206_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1206_/Y sky130_fd_sc_hd__inv_2
X_1068_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1068_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0918__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1331_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0706_ _0706_/A _0726_/A _0712_/A vssd1 vssd1 vccd1 vccd1 _0710_/A sky130_fd_sc_hd__and3_1
X_0637_ _0813_/A _0785_/A _0823_/A _0821_/A vssd1 vssd1 vccd1 vccd1 _0642_/D sky130_fd_sc_hd__or4bb_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0909__B2 hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 _0801_/X vssd1 vssd1 vccd1 vccd1 _1364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _0806_/X vssd1 vssd1 vccd1 vccd1 _1362_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _0808_/X vssd1 vssd1 vccd1 vccd1 _1361_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _0642_/C vssd1 vssd1 vccd1 vccd1 _0638_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _1355_/Q vssd1 vssd1 vccd1 vccd1 _0821_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold233 _1352_/Q vssd1 vssd1 vccd1 vccd1 _0785_/C sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold222 _1356_/Q vssd1 vssd1 vccd1 vccd1 _0813_/A sky130_fd_sc_hd__buf_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0898__B _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold288 _1400_/Q vssd1 vssd1 vccd1 vccd1 _0725_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _1399_/Q vssd1 vssd1 vccd1 vccd1 _0698_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _0735_/X vssd1 vssd1 vccd1 vccd1 _1396_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1014__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ hold14/X _0958_/X _0970_/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__a21o_1
X_1385_ _1386_/CLK hold43/X _1199_/Y vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1009__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1170_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1170_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0758__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0954_ hold163/X _0859_/D _0956_/S vssd1 vssd1 vccd1 vccd1 _1297_/D sky130_fd_sc_hd__mux2_1
X_0885_ _0875_/C _0884_/Y _0879_/D vssd1 vssd1 vccd1 vccd1 _0885_/X sky130_fd_sc_hd__a21o_1
X_1368_ _1419_/CLK _1368_/D _1182_/Y vssd1 vssd1 vccd1 vccd1 _1368_/Q sky130_fd_sc_hd__dfrtp_1
X_1299_ _1338_/CLK _1299_/D _1113_/Y vssd1 vssd1 vccd1 vccd1 _1299_/Q sky130_fd_sc_hd__dfrtp_1
Xinput15 wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_1
Xinput26 wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
X_0670_ _0749_/B _1408_/Q vssd1 vssd1 vccd1 vccd1 _0690_/A sky130_fd_sc_hd__nand2_1
X_1084_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1084_/Y sky130_fd_sc_hd__inv_2
X_1222_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1222_/Y sky130_fd_sc_hd__inv_2
X_1153_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1153_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0799_ _0802_/A _0802_/B vssd1 vssd1 vccd1 vccd1 _0799_/Y sky130_fd_sc_hd__nand2_1
X_0937_ hold115/X _0956_/S _0985_/B _1375_/Q vssd1 vssd1 vccd1 vccd1 _0937_/X sky130_fd_sc_hd__a22o_1
X_0868_ _1025_/A _1025_/C _0624_/Y vssd1 vssd1 vccd1 vccd1 _0868_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_3_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire94 wire94/A vssd1 vssd1 vccd1 vccd1 wire94/X sky130_fd_sc_hd__buf_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0653_ _0653_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0653_/X sky130_fd_sc_hd__or2_1
X_0722_ _1400_/Q _0724_/B _0715_/A vssd1 vssd1 vccd1 vccd1 _0722_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0945__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1136_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1136_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1067_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1067_/Y sky130_fd_sc_hd__inv_2
X_1205_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0936__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1017__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0636_ _0789_/A _0788_/A _0816_/S _1357_/Q vssd1 vssd1 vccd1 vccd1 _0642_/C sky130_fd_sc_hd__or4b_1
XANTENNA__0918__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0705_ _0673_/B _1405_/Q _0726_/A _0712_/A _0762_/S vssd1 vssd1 vccd1 vccd1 _0705_/Y
+ sky130_fd_sc_hd__a41oi_2
XFILLER_0_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1119_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1119_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0909__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold201 _1395_/Q vssd1 vssd1 vccd1 vccd1 _0693_/A sky130_fd_sc_hd__buf_1
Xhold234 _0828_/Y vssd1 vssd1 vccd1 vccd1 _0829_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _0822_/X vssd1 vssd1 vccd1 vccd1 _1355_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _0820_/X vssd1 vssd1 vccd1 vccd1 _1356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _1354_/Q vssd1 vssd1 vccd1 vccd1 _0785_/A sky130_fd_sc_hd__dlygate4sd3_1
X_0619_ _0647_/A vssd1 vssd1 vccd1 vccd1 _0653_/A sky130_fd_sc_hd__inv_2
Xhold289 _0725_/X vssd1 vssd1 vccd1 vccd1 _1400_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _0727_/X vssd1 vssd1 vccd1 vccd1 _0728_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _1398_/Q vssd1 vssd1 vccd1 vccd1 _0730_/A sky130_fd_sc_hd__buf_1
Xhold256 _1283_/Q vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0899__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1030__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1383_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0970_ _0958_/X hold97/A _0970_/C vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__and3b_1
X_1384_ _1390_/CLK hold88/X _1198_/Y vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0953_ _0864_/D _0853_/D _0956_/S vssd1 vssd1 vccd1 vccd1 _1298_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0884_ _0884_/A _0884_/B vssd1 vssd1 vccd1 vccd1 _0884_/Y sky130_fd_sc_hd__nand2_1
X_1367_ _1369_/CLK _1367_/D _1181_/Y vssd1 vssd1 vccd1 vccd1 _1367_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1298_ _1331_/CLK _1298_/D _1112_/Y vssd1 vssd1 vccd1 vccd1 _1298_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_1
XANTENNA__0957__A0 _0864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
X_1221_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1221_/Y sky130_fd_sc_hd__inv_2
X_1083_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1083_/Y sky130_fd_sc_hd__inv_2
X_1152_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1152_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0936_ hold73/X _0946_/A2 _0985_/B _1376_/Q vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__a22o_1
X_0798_ _0823_/D _0793_/Y _0797_/X _0796_/Y _0794_/A vssd1 vssd1 vccd1 vccd1 _0798_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout108_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0867_ _0850_/B _0866_/X _0867_/S vssd1 vssd1 vccd1 vccd1 _1347_/D sky130_fd_sc_hd__mux2_1
X_1419_ _1419_/CLK _1419_/D _1233_/Y vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0939__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0618__A hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0652_ _0652_/A hold57/X vssd1 vssd1 vccd1 vccd1 _0653_/B sky130_fd_sc_hd__nand2_1
X_0721_ _0723_/B _0720_/Y _0721_/S vssd1 vssd1 vccd1 vccd1 _0721_/X sky130_fd_sc_hd__mux2_1
X_1204_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1204_/Y sky130_fd_sc_hd__inv_2
X_1135_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1135_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1066_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1066_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0919_ _0931_/A _0919_/B vssd1 vssd1 vccd1 vccd1 _0919_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1033__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold172_A _1373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0635_ _0635_/A _0794_/A _0785_/C _1351_/Q vssd1 vssd1 vccd1 vccd1 _0642_/B sky130_fd_sc_hd__or4bb_1
X_0704_ _0726_/A _0704_/B vssd1 vssd1 vccd1 vccd1 _0733_/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1118_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1118_/Y sky130_fd_sc_hd__inv_2
X_1049_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1049_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1028__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold235 _0829_/Y vssd1 vssd1 vccd1 vccd1 _1352_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _0825_/X vssd1 vssd1 vccd1 vccd1 _1354_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold224 hold315/X vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__buf_1
Xhold202 _0737_/X vssd1 vssd1 vccd1 vccd1 _1395_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0618_ hold65/X vssd1 vssd1 vccd1 vccd1 _0891_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold279 _0728_/X vssd1 vssd1 vccd1 vccd1 _1399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _0731_/X vssd1 vssd1 vccd1 vccd1 _1398_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _1393_/Q vssd1 vssd1 vccd1 vccd1 _0742_/S sky130_fd_sc_hd__buf_1
Xhold257 _1236_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1383_ _1383_/CLK _1383_/D _1197_/Y vssd1 vssd1 vccd1 vccd1 _1383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0993__A1 _0864_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1041__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0952_ hold149/X _0860_/C _0956_/S vssd1 vssd1 vccd1 vccd1 _1299_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0975__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0883_ _0902_/B _0883_/B vssd1 vssd1 vccd1 vccd1 _0883_/X sky130_fd_sc_hd__and2_1
X_1366_ _1418_/CLK _1366_/D _1180_/Y vssd1 vssd1 vccd1 vccd1 _1366_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1297_ _1331_/CLK _1297_/D _1111_/Y vssd1 vssd1 vccd1 vccd1 _1297_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0966__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1386_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__1036__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
Xinput28 wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
X_1151_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1151_/Y sky130_fd_sc_hd__inv_2
X_1220_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1220_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0893__B1 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1082_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1082_/Y sky130_fd_sc_hd__inv_2
X_0935_ hold145/X _0948_/A2 _0985_/B _1377_/Q vssd1 vssd1 vccd1 vccd1 _0935_/X sky130_fd_sc_hd__a22o_1
X_0866_ hold149/X hold55/X hold186/X _0865_/X _0861_/X vssd1 vssd1 vccd1 vccd1 _0866_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0797_ _0794_/C _0802_/B _0794_/A vssd1 vssd1 vccd1 vccd1 _0797_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1418_ _1418_/CLK _1418_/D _1232_/Y vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfrtp_1
X_1349_ _1407_/CLK input2/X _1163_/Y vssd1 vssd1 vccd1 vccd1 _1349_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__0724__A _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0939__B2 _1373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0720_ _0720_/A _0720_/B vssd1 vssd1 vccd1 vccd1 _0720_/Y sky130_fd_sc_hd__nor2_1
X_0651_ _0656_/A _0651_/B vssd1 vssd1 vccd1 vccd1 _0651_/Y sky130_fd_sc_hd__nor2_1
X_1134_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1134_/Y sky130_fd_sc_hd__inv_2
X_1203_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1203_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1065_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1065_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0918_ hold147/X _0948_/A2 _0917_/Y _0908_/B vssd1 vssd1 vccd1 vccd1 _0918_/X sky130_fd_sc_hd__a22o_1
X_0849_ _0849_/A _0849_/B _0852_/B vssd1 vssd1 vccd1 vccd1 _0892_/B sky130_fd_sc_hd__nor3_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0703_ _0726_/A _0704_/B vssd1 vssd1 vccd1 vccd1 _0762_/S sky130_fd_sc_hd__nor2_8
X_0634_ _0784_/A _0791_/A _0807_/A _0802_/A vssd1 vssd1 vccd1 vccd1 _0642_/A sky130_fd_sc_hd__or4bb_1
X_1117_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1117_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1048_ _1048_/A _1048_/B vssd1 vssd1 vccd1 vccd1 _1390_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold258 hold314/X vssd1 vssd1 vccd1 vccd1 _0802_/A sky130_fd_sc_hd__buf_1
Xhold236 _1366_/Q vssd1 vssd1 vccd1 vccd1 _0635_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _1358_/Q vssd1 vssd1 vccd1 vccd1 _0816_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold203 _1319_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _1284_/Q vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _1018_/X vssd1 vssd1 vccd1 vccd1 _1256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _0742_/X vssd1 vssd1 vccd1 vccd1 _1393_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0617_ _0700_/A vssd1 vssd1 vccd1 vccd1 _0717_/A sky130_fd_sc_hd__inv_2
XANTENNA__1039__S _1041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1382_ _1411_/CLK hold21/X _1196_/Y vssd1 vssd1 vccd1 vccd1 _1382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0951_ _0863_/B _0853_/B _0956_/S vssd1 vssd1 vccd1 vccd1 _1300_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0882_ _0875_/X _0882_/B _0882_/C vssd1 vssd1 vccd1 vccd1 _1344_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1365_ _1418_/CLK _1365_/D _1179_/Y vssd1 vssd1 vccd1 vccd1 _1365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1296_ _1331_/CLK _1296_/D _1110_/Y vssd1 vssd1 vccd1 vccd1 _1296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
Xinput29 wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
X_1150_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1150_/Y sky130_fd_sc_hd__inv_2
X_1081_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1081_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0948__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0865_ _0891_/A _0863_/B _0864_/X _0863_/Y vssd1 vssd1 vccd1 vccd1 _0865_/X sky130_fd_sc_hd__a31o_1
X_0934_ hold61/X _0946_/A2 _0985_/B hold65/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__a22o_1
X_0796_ input1/X _0813_/C vssd1 vssd1 vccd1 vccd1 _0796_/Y sky130_fd_sc_hd__nor2_2
X_1417_ _1417_/CLK hold60/X _1231_/Y vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1348_ _1348_/CLK _1348_/D _1162_/Y vssd1 vssd1 vccd1 vccd1 _1348_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1279_ _1404_/CLK _1279_/D _1093_/Y vssd1 vssd1 vccd1 vccd1 _1279_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0939__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold208_A _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0897__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0650_ _0629_/Y hold49/X _0649_/Y _0644_/X vssd1 vssd1 vccd1 vccd1 _1419_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1133_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1133_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0866__A1 hold149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1202_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1202_/Y sky130_fd_sc_hd__inv_2
X_1064_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1064_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1338_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0917_ _0931_/A hold92/X vssd1 vssd1 vccd1 vccd1 _0917_/Y sky130_fd_sc_hd__nor2_1
X_0779_ _0640_/B _0775_/Y _0764_/B _0653_/B vssd1 vssd1 vccd1 vccd1 _0779_/Y sky130_fd_sc_hd__a211oi_1
X_0848_ _0884_/A _0933_/B _0846_/X _0847_/X vssd1 vssd1 vccd1 vccd1 _1025_/C sky130_fd_sc_hd__a211oi_2
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0633_ _0647_/A _0632_/A hold79/X vssd1 vssd1 vccd1 vccd1 _0763_/B sky130_fd_sc_hd__o21a_1
X_0702_ _1406_/Q _1405_/Q _0726_/A _0712_/A vssd1 vssd1 vccd1 vccd1 _0702_/X sky130_fd_sc_hd__and4_1
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1116_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1116_/Y sky130_fd_sc_hd__inv_2
X_1047_ _0813_/C _1046_/X _0773_/S vssd1 vssd1 vccd1 vccd1 _1350_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold237 _0642_/B vssd1 vssd1 vccd1 vccd1 _0638_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _0816_/X vssd1 vssd1 vccd1 vccd1 _1358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _1353_/Q vssd1 vssd1 vccd1 vccd1 _0823_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _1020_/X vssd1 vssd1 vccd1 vccd1 _1254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 _1279_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold248 _1394_/Q vssd1 vssd1 vccd1 vccd1 _0740_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0911__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1381_ _1411_/CLK hold45/X _1195_/Y vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0978__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0950_ hold65/X _0860_/D _0956_/S vssd1 vssd1 vccd1 vccd1 _1301_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0881_ _0883_/B _0879_/D hold96/X vssd1 vssd1 vccd1 vccd1 _0882_/C sky130_fd_sc_hd__a21o_1
X_1364_ _1418_/CLK _1364_/D _1178_/Y vssd1 vssd1 vccd1 vccd1 _1364_/Q sky130_fd_sc_hd__dfrtp_1
X_1295_ _1331_/CLK _1295_/D _1109_/Y vssd1 vssd1 vccd1 vccd1 _1295_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
X_1080_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1080_/Y sky130_fd_sc_hd__inv_2
X_0795_ _0783_/Y _0783_/A _0795_/S vssd1 vssd1 vccd1 vccd1 _1366_/D sky130_fd_sc_hd__mux2_1
X_0864_ _1374_/Q _0864_/B _0864_/C _0864_/D vssd1 vssd1 vccd1 vccd1 _0864_/X sky130_fd_sc_hd__and4b_1
X_0933_ _0884_/A _0933_/B vssd1 vssd1 vccd1 vccd1 _0985_/B sky130_fd_sc_hd__and2b_4
X_1416_ _1419_/CLK _1416_/D _1230_/Y vssd1 vssd1 vccd1 vccd1 _1416_/Q sky130_fd_sc_hd__dfrtp_1
X_1347_ _1348_/CLK _1347_/D _1161_/Y vssd1 vssd1 vccd1 vccd1 _1347_/Q sky130_fd_sc_hd__dfrtp_1
X_1278_ _1418_/CLK _1278_/D _1092_/Y vssd1 vssd1 vccd1 vccd1 _1278_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0992__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1201_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1201_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1132_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1132_/Y sky130_fd_sc_hd__inv_2
X_1063_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1063_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0866__A2 hold55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0916_ hold138/X _0946_/A2 _0908_/X _0864_/C vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0778_ hold79/X _0777_/X _0655_/S vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout106_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0847_ _0892_/A _1025_/B vssd1 vssd1 vccd1 vccd1 _0847_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0632_ _0632_/A _0668_/A vssd1 vssd1 vccd1 vccd1 _0643_/A sky130_fd_sc_hd__nor2_1
X_0701_ _0701_/A _0719_/B _0701_/C vssd1 vssd1 vccd1 vccd1 _0712_/A sky130_fd_sc_hd__and3_1
XFILLER_0_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1046_ hold48/X input1/X vssd1 vssd1 vccd1 vccd1 _1046_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1115_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1115_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0766__A1 hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1339_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold205 _1257_/Q vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 _1303_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _0642_/X vssd1 vssd1 vccd1 vccd1 _0803_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _0827_/X vssd1 vssd1 vccd1 vccd1 _1353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _0740_/X vssd1 vssd1 vccd1 vccd1 _1394_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0996__A1 hold55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1029_ hold124/X hold115/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1029_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0920__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1380_ _1390_/CLK _1380_/D _1194_/Y vssd1 vssd1 vccd1 vccd1 _1380_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0911__B2 hold149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0995__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0969__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0880_ _0878_/X _0879_/Y _0875_/X vssd1 vssd1 vccd1 vccd1 _1345_/D sky130_fd_sc_hd__a21oi_1
X_1363_ _1369_/CLK _1363_/D _1177_/Y vssd1 vssd1 vccd1 vccd1 _1363_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1294_ _1348_/CLK _1294_/D _1108_/Y vssd1 vssd1 vccd1 vccd1 _1294_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0887__B1 _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0932_ hold119/X _0956_/S _0931_/Y _0908_/B vssd1 vssd1 vccd1 vccd1 _0932_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0794_ _0794_/A _0823_/D _0794_/C _0802_/B vssd1 vssd1 vccd1 vccd1 _0795_/S sky130_fd_sc_hd__and4_1
X_0863_ _0891_/A _0863_/B _0863_/C vssd1 vssd1 vccd1 vccd1 _0863_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1415_ _1417_/CLK _1415_/D _1229_/Y vssd1 vssd1 vccd1 vccd1 _1415_/Q sky130_fd_sc_hd__dfrtp_1
X_1346_ _1348_/CLK _1346_/D _1160_/Y vssd1 vssd1 vccd1 vccd1 _1346_/Q sky130_fd_sc_hd__dfrtp_1
X_1277_ _1386_/CLK _1277_/D _1091_/Y vssd1 vssd1 vccd1 vccd1 _1277_/Q sky130_fd_sc_hd__dfrtp_1
X_1200_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1200_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1131_/Y sky130_fd_sc_hd__inv_2
X_1062_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1062_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0915_ hold2/X _0946_/A2 _0908_/X hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__a22o_1
X_0777_ _0823_/D _0654_/B _0775_/Y _0640_/B _0764_/B vssd1 vssd1 vccd1 vccd1 _0777_/X
+ sky130_fd_sc_hd__a221o_1
X_0846_ hold96/X _0890_/B _0989_/A _0889_/B vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__o31a_1
X_1329_ _1338_/CLK hold39/X _1143_/Y vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ _0700_/A _0721_/S _0715_/A _1400_/Q vssd1 vssd1 vccd1 vccd1 _0701_/C sky130_fd_sc_hd__and4_1
X_0631_ hold79/X _0647_/A vssd1 vssd1 vccd1 vccd1 _0668_/A sky130_fd_sc_hd__or2_2
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1114_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1114_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1045_ _0835_/B _0733_/A _1048_/B vssd1 vssd1 vccd1 vccd1 _1045_/X sky130_fd_sc_hd__a21o_1
XANTENNA__0998__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0829_ _0829_/A _0829_/B vssd1 vssd1 vccd1 vccd1 _0829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold163_A _1374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 _1348_/Q vssd1 vssd1 vccd1 vccd1 _0852_/C sky130_fd_sc_hd__buf_2
Xhold217 _1404_/Q vssd1 vssd1 vccd1 vccd1 _0701_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold239 _0668_/B vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _1343_/Q vssd1 vssd1 vccd1 vccd1 _0841_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1028_ hold100/X hold73/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0895__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1362_ _1369_/CLK _1362_/D _1176_/Y vssd1 vssd1 vccd1 vccd1 _1362_/Q sky130_fd_sc_hd__dfrtp_1
X_1293_ _1411_/CLK hold17/X _1107_/Y vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0754__B _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0931_ _0931_/A _0931_/B vssd1 vssd1 vccd1 vccd1 _0931_/Y sky130_fd_sc_hd__nor2_1
X_0862_ _1375_/Q _1373_/Q _1371_/Q _1374_/Q vssd1 vssd1 vccd1 vccd1 _0863_/C sky130_fd_sc_hd__or4b_1
X_0793_ _0794_/A _0794_/C _0802_/B vssd1 vssd1 vccd1 vccd1 _0793_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1276_ _1341_/CLK hold86/X _1090_/Y vssd1 vssd1 vccd1 vccd1 _1276_/Q sky130_fd_sc_hd__dfrtp_2
X_1414_ _1419_/CLK _1414_/D _1228_/Y vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfrtp_1
X_1345_ _1383_/CLK _1345_/D _1159_/Y vssd1 vssd1 vccd1 vccd1 _1345_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0839__B _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout110 input3/X vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1130_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1130_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1061_ _1139_/A vssd1 vssd1 vccd1 vccd1 _1061_/Y sky130_fd_sc_hd__inv_2
X_0914_ hold71/X _0946_/A2 _0908_/X _0864_/B vssd1 vssd1 vccd1 vccd1 _0914_/X sky130_fd_sc_hd__a22o_1
X_0845_ _0852_/C _0850_/B _0852_/B vssd1 vssd1 vccd1 vccd1 _0889_/B sky130_fd_sc_hd__and3b_2
X_0776_ _0640_/B _0775_/Y _0764_/B vssd1 vssd1 vccd1 vccd1 _0776_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1259_ _1340_/CLK _1259_/D _1073_/Y vssd1 vssd1 vccd1 vccd1 _1259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1328_ _1411_/CLK _1328_/D _1142_/Y vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0950__A0 hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0941__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0630_ _0652_/A hold57/X vssd1 vssd1 vccd1 vccd1 _0632_/A sky130_fd_sc_hd__or2_2
X_1044_ _0749_/A _0749_/B _0726_/A _0678_/C _0745_/A vssd1 vssd1 vccd1 vccd1 _1048_/B
+ sky130_fd_sc_hd__o2111a_1
X_1113_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1113_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0828_ _1351_/Q _0823_/D _0785_/C vssd1 vssd1 vccd1 vccd1 _0828_/Y sky130_fd_sc_hd__a21oi_1
X_0759_ hold106/X hold10/X _0762_/S vssd1 vssd1 vccd1 vccd1 _0759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold229 hold312/X vssd1 vssd1 vccd1 vccd1 _0652_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 _0713_/X vssd1 vssd1 vccd1 vccd1 _1404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold207 _0889_/B vssd1 vssd1 vccd1 vccd1 _0857_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0914__B1 _0908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1027_ hold164/X hold145/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1251_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0905__B1 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout91_A _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1361_ _1369_/CLK _1361_/D _1175_/Y vssd1 vssd1 vccd1 vccd1 _1361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1292_ _1386_/CLK hold7/X _1106_/Y vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfrtp_1
Xoutput80 _1256_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[3] sky130_fd_sc_hd__buf_12
XANTENNA__0902__C_N _1373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0792_ _0794_/C _0802_/B vssd1 vssd1 vccd1 vccd1 _0792_/Y sky130_fd_sc_hd__nand2_1
X_0930_ hold203/X _0956_/S _0929_/Y hold208/X vssd1 vssd1 vccd1 vccd1 _1319_/D sky130_fd_sc_hd__a22o_1
X_0861_ _0884_/B _0859_/X _0860_/X _0871_/D vssd1 vssd1 vccd1 vccd1 _0861_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1413_ _1419_/CLK _1413_/D _1227_/Y vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfrtp_1
X_1275_ _1341_/CLK _1275_/D _1089_/Y vssd1 vssd1 vccd1 vccd1 _1275_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1344_ _1383_/CLK _1344_/D _1158_/Y vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout111 _1233_/A vssd1 vssd1 vccd1 vccd1 _1232_/A sky130_fd_sc_hd__buf_8
Xfanout100 _1197_/A vssd1 vssd1 vccd1 vccd1 _1153_/A sky130_fd_sc_hd__buf_8
X_1060_ _1231_/A vssd1 vssd1 vccd1 vccd1 _1060_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0775_ _0813_/C input1/X vssd1 vssd1 vccd1 vccd1 _0775_/Y sky130_fd_sc_hd__nand2b_1
X_0844_ _0852_/C _0850_/B vssd1 vssd1 vccd1 vccd1 _1025_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0913_ hold38/X _0946_/A2 _0908_/X _1374_/Q vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__a22o_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1258_ _1418_/CLK hold47/X _1072_/Y vssd1 vssd1 vccd1 vccd1 _1258_/Q sky130_fd_sc_hd__dfrtp_2
X_1189_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1189_/Y sky130_fd_sc_hd__inv_2
X_1327_ _1338_/CLK hold56/X _1141_/Y vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0769__A1 _1375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0941__B2 _0864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1043_ hold303/X _1025_/B _1043_/S vssd1 vssd1 vccd1 vccd1 _1235_/D sky130_fd_sc_hd__mux2_1
X_1112_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1112_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ _0823_/A _0829_/A _0823_/X vssd1 vssd1 vccd1 vccd1 _0827_/X sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout104_A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0758_ hold87/X hold14/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__mux2_1
XANTENNA__0932__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0689_ _0749_/B _1408_/Q vssd1 vssd1 vccd1 vccd1 _0690_/B sky130_fd_sc_hd__or2_1
Xhold208 _0908_/B vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold219 _1406_/Q vssd1 vssd1 vccd1 vccd1 _0673_/B sky130_fd_sc_hd__buf_1
XFILLER_0_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0914__B2 _0864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1026_ _1252_/Q hold61/X _1041_/S vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__mux2_1
XFILLER_0_31_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0899__B1 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1009_ hold165/X hold128/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1265_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput70 _1276_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[23] sky130_fd_sc_hd__buf_12
X_1360_ _1369_/CLK _1360_/D _1174_/Y vssd1 vssd1 vccd1 vccd1 _1360_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput81 _1257_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[4] sky130_fd_sc_hd__buf_12
X_1291_ _1383_/CLK hold27/X _1105_/Y vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfrtp_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0791_ _0791_/A _0807_/A _0807_/B vssd1 vssd1 vccd1 vccd1 _0802_/B sky130_fd_sc_hd__and3_2
X_0860_ _0853_/B _0853_/D _0860_/C _0860_/D vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_48_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1412_ _1417_/CLK hold50/X _1226_/Y vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfrtp_1
X_1343_ _1383_/CLK _1343_/D _1157_/Y vssd1 vssd1 vccd1 vccd1 _1343_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1274_ _1339_/CLK _1274_/D _1088_/Y vssd1 vssd1 vccd1 vccd1 _1274_/Q sky130_fd_sc_hd__dfrtp_1
X_0989_ _0989_/A _0989_/B vssd1 vssd1 vccd1 vccd1 _1003_/S sky130_fd_sc_hd__nor2_2
Xfanout112 _1233_/A vssd1 vssd1 vccd1 vccd1 _1180_/A sky130_fd_sc_hd__buf_8
Xfanout101 _1197_/A vssd1 vssd1 vccd1 vccd1 _1158_/A sky130_fd_sc_hd__buf_8
XFILLER_0_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0907__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0912_ hold128/X _0956_/S _0908_/X _1375_/Q vssd1 vssd1 vccd1 vccd1 _0912_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0774_ _0813_/C input1/X vssd1 vssd1 vccd1 vccd1 _0815_/A sky130_fd_sc_hd__and2b_2
X_0843_ _0849_/A hold309/X _0892_/A _0849_/B vssd1 vssd1 vccd1 vccd1 _0933_/B sky130_fd_sc_hd__and4bb_4
X_1326_ _1411_/CLK _1326_/D _1140_/Y vssd1 vssd1 vccd1 vccd1 _1326_/Q sky130_fd_sc_hd__dfrtp_1
X_1257_ _1341_/CLK _1257_/D _1071_/Y vssd1 vssd1 vccd1 vccd1 _1257_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0893__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1188_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1188_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0941__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1111_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1111_/Y sky130_fd_sc_hd__inv_2
X_1042_ hold257/X _0857_/A _1042_/S vssd1 vssd1 vccd1 vccd1 _1236_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0826_ _0785_/C _1351_/Q _0823_/D _0815_/A vssd1 vssd1 vccd1 vccd1 _0829_/A sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_4_6_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0757_ hold42/X hold26/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__mux2_1
X_0688_ _0749_/A _0685_/Y _0687_/X vssd1 vssd1 vccd1 vccd1 _0688_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_4_15_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1369_/CLK sky130_fd_sc_hd__clkbuf_8
X_1309_ _1331_/CLK _1309_/D _1123_/Y vssd1 vssd1 vccd1 vccd1 _1309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold209 _1295_/Q vssd1 vssd1 vccd1 vccd1 _0859_/C sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0914__A2 _0946_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1025_ _1025_/A _1025_/B _1025_/C _1025_/D vssd1 vssd1 vccd1 vccd1 _1041_/S sky130_fd_sc_hd__and4_4
X_0809_ input1/X _0788_/X _0813_/C vssd1 vssd1 vccd1 vccd1 _0809_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold161_A _1343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _1266_/Q hold176/X _1021_/S vssd1 vssd1 vccd1 vccd1 _1008_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput82 _1258_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[5] sky130_fd_sc_hd__buf_12
Xoutput71 _1277_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput60 _1267_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[14] sky130_fd_sc_hd__buf_12
X_1290_ _1390_/CLK hold15/X _1104_/Y vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0790_ _0807_/A _0807_/B vssd1 vssd1 vccd1 vccd1 _0790_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1411_ _1411_/CLK _1411_/D _1225_/Y vssd1 vssd1 vccd1 vccd1 _1411_/Q sky130_fd_sc_hd__dfrtp_1
X_1273_ _1339_/CLK hold5/X _1087_/Y vssd1 vssd1 vccd1 vccd1 _1273_/Q sky130_fd_sc_hd__dfrtp_2
X_1342_ _1383_/CLK _1342_/D _1156_/Y vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0988_ _1025_/C _0988_/B _0988_/C _0988_/D vssd1 vssd1 vccd1 vccd1 _1042_/S sky130_fd_sc_hd__and4_1
Xfanout113 _1233_/A vssd1 vssd1 vccd1 vccd1 _1178_/A sky130_fd_sc_hd__buf_4
Xfanout102 _1197_/A vssd1 vssd1 vccd1 vccd1 _1225_/A sky130_fd_sc_hd__buf_8
XANTENNA__0953__A0 _0864_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0705__B1 _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0862__D_N _1374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0911_ hold176/X _0956_/S _0908_/X hold149/X vssd1 vssd1 vccd1 vccd1 _1331_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0842_ _0852_/C _0871_/A vssd1 vssd1 vccd1 vccd1 _0884_/B sky130_fd_sc_hd__and2b_1
X_0773_ hold34/X _1371_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__mux2_1
X_1325_ _1340_/CLK _1325_/D _1139_/Y vssd1 vssd1 vccd1 vccd1 _1325_/Q sky130_fd_sc_hd__dfrtp_1
X_1256_ _1383_/CLK _1256_/D _1070_/Y vssd1 vssd1 vccd1 vccd1 _1256_/Q sky130_fd_sc_hd__dfrtp_1
X_1187_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1187_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_2_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0935__B1 _0985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1162_/A vssd1 vssd1 vccd1 vccd1 _1110_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1041_ hold122/X hold94/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1041_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0825_ _0785_/A _0815_/A _0823_/X _0824_/Y vssd1 vssd1 vccd1 vccd1 _0825_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0756_ hold40/X hold6/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0687_ _0749_/A _0690_/A _0687_/C vssd1 vssd1 vccd1 vccd1 _0687_/X sky130_fd_sc_hd__or3_1
X_1308_ _1340_/CLK _1308_/D _1122_/Y vssd1 vssd1 vccd1 vccd1 _1308_/Q sky130_fd_sc_hd__dfrtp_1
X_1239_ _1340_/CLK _1239_/D _1053_/Y vssd1 vssd1 vccd1 vccd1 _1239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1024_ _1025_/A _1025_/C _1025_/D vssd1 vssd1 vccd1 vccd1 _1043_/S sky130_fd_sc_hd__and3_1
XFILLER_0_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0808_ _0790_/Y _0803_/X _0807_/X _0796_/Y _0807_/A vssd1 vssd1 vccd1 vccd1 _0808_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0739_ _0762_/S _0739_/B vssd1 vssd1 vccd1 vccd1 _0739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1419_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0864__A_N _1374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1007_ hold110/X hold63/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1267_/D sky130_fd_sc_hd__mux2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput83 _1259_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xoutput72 _1278_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput50 _1243_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[6] sky130_fd_sc_hd__buf_12
Xoutput61 _1268_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1001__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1410_ _1411_/CLK _1410_/D _1224_/Y vssd1 vssd1 vccd1 vccd1 _1410_/Q sky130_fd_sc_hd__dfrtp_1
X_1272_ _1341_/CLK _1272_/D _1086_/Y vssd1 vssd1 vccd1 vccd1 _1272_/Q sky130_fd_sc_hd__dfrtp_2
X_1341_ _1341_/CLK hold93/X _1155_/Y vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0987_ _0850_/B _0892_/A _0624_/Y _0852_/C vssd1 vssd1 vccd1 vccd1 _0988_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout114 input3/X vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout103 _1197_/A vssd1 vssd1 vccd1 vccd1 _1218_/A sky130_fd_sc_hd__buf_4
Xhold190 _1296_/Q vssd1 vssd1 vccd1 vccd1 _0854_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0772_ hold18/X _1372_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__mux2_1
X_0910_ hold63/X _0946_/A2 _0908_/X _1377_/Q vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__a22o_1
X_0841_ _0906_/A hold96/X _0841_/C _0902_/B vssd1 vssd1 vccd1 vccd1 _0884_/A sky130_fd_sc_hd__or4b_2
X_1324_ _1340_/CLK _1324_/D _1138_/Y vssd1 vssd1 vccd1 vccd1 _1324_/Q sky130_fd_sc_hd__dfrtp_1
X_1186_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1186_/Y sky130_fd_sc_hd__inv_2
X_1255_ _1339_/CLK _1255_/D _1069_/Y vssd1 vssd1 vccd1 vccd1 _1255_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0935__B2 _1377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0926__B2 _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1040_ hold221/X hold216/X _1041_/S vssd1 vssd1 vccd1 vccd1 _1238_/D sky130_fd_sc_hd__mux2_1
X_0824_ _0638_/Y _0821_/B _0823_/D vssd1 vssd1 vccd1 vccd1 _0824_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0755_ hold28/X hold16/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__mux2_1
XFILLER_0_9_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0686_ _0678_/X _0685_/Y _0745_/A vssd1 vssd1 vccd1 vccd1 _0686_/X sky130_fd_sc_hd__mux2_1
X_1169_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1169_/Y sky130_fd_sc_hd__inv_2
X_1307_ _1341_/CLK _1307_/D _1121_/Y vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfrtp_1
X_1238_ _1418_/CLK _1238_/D _1052_/Y vssd1 vssd1 vccd1 vccd1 _1238_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1023_ _0985_/A _0985_/B _1022_/X vssd1 vssd1 vccd1 vccd1 _1025_/D sky130_fd_sc_hd__a21boi_1
X_0807_ _0807_/A _0807_/B vssd1 vssd1 vccd1 vccd1 _0807_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout102_A _1197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0738_ _0742_/S _1392_/Q _1390_/Q vssd1 vssd1 vccd1 vccd1 _0739_/B sky130_fd_sc_hd__and3_1
X_0669_ hold49/X hold34/X _0669_/S vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
XANTENNA__1004__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0905__A1_N _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ hold132/X hold104/X _1019_/S vssd1 vssd1 vccd1 vccd1 _1268_/D sky130_fd_sc_hd__mux2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput84 _1260_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[7] sky130_fd_sc_hd__buf_12
Xoutput73 _1279_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput62 _1269_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput40 hold83/A vssd1 vssd1 vccd1 vccd1 wb_adr_o[11] sky130_fd_sc_hd__buf_12
Xoutput51 _1244_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1418_/CLK sky130_fd_sc_hd__clkbuf_8
X_1340_ _1340_/CLK _1340_/D _1154_/Y vssd1 vssd1 vccd1 vccd1 _1340_/Q sky130_fd_sc_hd__dfrtp_1
X_1271_ _1341_/CLK _1271_/D _1085_/Y vssd1 vssd1 vccd1 vccd1 _1271_/Q sky130_fd_sc_hd__dfrtp_1
X_0986_ _0850_/B _0837_/B _0852_/C vssd1 vssd1 vccd1 vccd1 _0988_/C sky130_fd_sc_hd__o21ai_1
Xfanout104 _1197_/A vssd1 vssd1 vccd1 vccd1 _1231_/A sky130_fd_sc_hd__buf_8
XANTENNA__0896__B _0902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1012__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 _1339_/Q vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0890__C_N _0908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 _1298_/Q vssd1 vssd1 vccd1 vccd1 _0853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0771_ hold69/X _1373_/Q _0773_/S vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__mux2_1
XANTENNA__0761__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0840_ hold96/X _0876_/A vssd1 vssd1 vccd1 vccd1 _0931_/A sky130_fd_sc_hd__or2_4
X_1323_ _1341_/CLK _1323_/D _1137_/Y vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__0944__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1254_ _1331_/CLK _1254_/D _1068_/Y vssd1 vssd1 vccd1 vccd1 _1254_/Q sky130_fd_sc_hd__dfrtp_1
X_1185_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1185_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0935__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0969_ input31/X input8/X input17/X input25/X hold91/A _1343_/Q vssd1 vssd1 vccd1
+ vccd1 _0970_/C sky130_fd_sc_hd__mux4_1
XANTENNA__1007__S _1019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0926__A2 _0948_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0756__S _0762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0823_ _0823_/A _1352_/Q _1351_/Q _0823_/D vssd1 vssd1 vccd1 vccd1 _0823_/X sky130_fd_sc_hd__and4_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0754_ hold8/X _0762_/S vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__or2_1
X_0685_ _0678_/B _0687_/C _0720_/A vssd1 vssd1 vccd1 vccd1 _0685_/Y sky130_fd_sc_hd__o21ai_1
X_1306_ _1338_/CLK hold76/X _1120_/Y vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfrtp_1
X_1168_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1168_/Y sky130_fd_sc_hd__inv_2
X_1237_ _1348_/CLK _1237_/D _1051_/Y vssd1 vssd1 vccd1 vccd1 _1237_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1099_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1099_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1022_ _0884_/A _0933_/B _1025_/B _0624_/Y vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0806_ _0823_/D _0802_/B _0805_/X _0791_/A vssd1 vssd1 vccd1 vccd1 _0806_/X sky130_fd_sc_hd__o2bb2a_1
X_0668_ _0668_/A _0668_/B _0645_/Y vssd1 vssd1 vccd1 vccd1 _0669_/S sky130_fd_sc_hd__or3b_1
X_0737_ _0684_/B _0694_/Y _0736_/X _1048_/A _0693_/A vssd1 vssd1 vccd1 vccd1 _0737_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1020__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0989__B _0989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _1269_/Q hold12/X _1019_/S vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1015__S _1021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput52 _1245_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[8] sky130_fd_sc_hd__buf_12
Xoutput41 _1249_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[12] sky130_fd_sc_hd__buf_12
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput63 _1270_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[17] sky130_fd_sc_hd__buf_12
Xoutput74 _1280_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput85 _1261_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[8] sky130_fd_sc_hd__buf_12
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

