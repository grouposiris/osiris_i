VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO osiris_i_mem
  CLASS BLOCK ;
  FOREIGN osiris_i_mem ;
  ORIGIN 0.000 0.000 ;
  SIZE 1356.000 BY 1120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1352.000 608.640 1356.000 609.240 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 550.710 1116.000 550.990 1120.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 872.710 1116.000 872.990 1120.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_in[4]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1352.000 948.640 1356.000 949.240 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 1116.000 1194.990 1120.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END io_oeb[6]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 1116.000 228.990 1120.000 ;
    END
  END io_out[1]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.200 6.000 30.800 1114.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 29.200 6.000 1340.220 7.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 29.200 1113.040 1340.220 1114.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.620 6.000 1340.220 1114.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.320 2.700 53.920 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 205.920 2.700 207.520 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 205.920 526.520 207.520 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 205.920 1042.520 207.520 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.520 2.700 361.120 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.520 526.520 361.120 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.520 1042.520 361.120 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.120 2.700 514.720 89.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.120 527.140 514.720 605.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.120 1043.140 514.720 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.720 2.700 668.320 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.720 527.140 668.320 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.720 1043.140 668.320 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 820.320 2.700 821.920 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 973.920 2.700 975.520 371.375 ;
    END
    PORT
      LAYER met4 ;
        RECT 973.920 1017.145 975.520 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1127.520 2.700 1129.120 371.375 ;
    END
    PORT
      LAYER met4 ;
        RECT 1127.520 1017.145 1129.120 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.120 2.700 1282.720 1117.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 29.450 1343.520 31.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 182.630 1343.520 184.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 335.810 1343.520 337.410 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 488.990 1343.520 490.590 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 642.170 1343.520 643.770 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 795.350 1343.520 796.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 948.530 1343.520 950.130 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 1101.710 1343.520 1103.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 1310.660 356.080 1312.260 1036.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 52.320 565.300 825.220 566.900 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.900 2.700 27.500 1117.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 2.700 1343.520 4.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 1116.340 1343.520 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1341.920 2.700 1343.520 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.620 2.700 57.220 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.220 2.700 210.820 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.220 526.520 210.820 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.220 1042.520 210.820 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 362.820 2.700 364.420 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 362.820 526.520 364.420 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 362.820 1042.520 364.420 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.420 2.700 518.020 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.420 527.140 518.020 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.420 1043.140 518.020 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 670.020 2.700 671.620 90.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 670.020 526.520 671.620 606.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 670.020 1042.520 671.620 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.620 2.700 825.220 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 977.220 2.700 978.820 371.375 ;
    END
    PORT
      LAYER met4 ;
        RECT 977.220 1017.145 978.820 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1130.820 2.700 1132.420 371.375 ;
    END
    PORT
      LAYER met4 ;
        RECT 1130.820 1017.145 1132.420 1117.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1284.420 2.700 1286.020 1117.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 32.750 1343.520 34.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 185.930 1343.520 187.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 339.110 1343.520 340.710 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 492.290 1343.520 493.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 645.470 1343.520 647.070 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 798.650 1343.520 800.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 951.830 1343.520 953.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.900 1105.010 1343.520 1106.610 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.340 356.080 1315.940 1036.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 52.320 568.700 825.220 570.300 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1352.000 268.640 1356.000 269.240 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 36.800 13.515 1332.620 1107.125 ;
      LAYER met1 ;
        RECT 0.070 13.360 1334.850 1107.280 ;
      LAYER met2 ;
        RECT 0.100 1115.720 228.430 1116.000 ;
        RECT 229.270 1115.720 550.430 1116.000 ;
        RECT 551.270 1115.720 872.430 1116.000 ;
        RECT 873.270 1115.720 1194.430 1116.000 ;
        RECT 1195.270 1115.720 1335.290 1116.000 ;
        RECT 0.100 4.280 1335.290 1115.720 ;
        RECT 0.650 4.000 321.810 4.280 ;
        RECT 322.650 4.000 643.810 4.280 ;
        RECT 644.650 4.000 965.810 4.280 ;
        RECT 966.650 4.000 1291.030 4.280 ;
        RECT 1291.870 4.000 1335.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 1021.040 1352.000 1107.205 ;
        RECT 4.400 1019.640 1352.000 1021.040 ;
        RECT 4.000 949.640 1352.000 1019.640 ;
        RECT 4.000 948.240 1351.600 949.640 ;
        RECT 4.000 681.040 1352.000 948.240 ;
        RECT 4.400 679.640 1352.000 681.040 ;
        RECT 4.000 609.640 1352.000 679.640 ;
        RECT 4.000 608.240 1351.600 609.640 ;
        RECT 4.000 341.040 1352.000 608.240 ;
        RECT 4.400 339.640 1352.000 341.040 ;
        RECT 4.000 269.640 1352.000 339.640 ;
        RECT 4.000 268.240 1351.600 269.640 ;
        RECT 4.000 13.435 1352.000 268.240 ;
      LAYER met4 ;
        RECT 100.620 1042.120 205.520 1105.505 ;
        RECT 207.920 1042.120 208.820 1105.505 ;
        RECT 211.220 1042.120 359.120 1105.505 ;
        RECT 361.520 1042.120 362.420 1105.505 ;
        RECT 364.820 1042.740 512.720 1105.505 ;
        RECT 515.120 1042.740 516.020 1105.505 ;
        RECT 518.420 1042.740 666.320 1105.505 ;
        RECT 668.720 1042.740 669.620 1105.505 ;
        RECT 364.820 1042.120 669.620 1042.740 ;
        RECT 672.020 1042.120 819.920 1105.505 ;
        RECT 100.620 606.420 819.920 1042.120 ;
        RECT 100.620 526.120 205.520 606.420 ;
        RECT 207.920 526.120 208.820 606.420 ;
        RECT 211.220 526.120 359.120 606.420 ;
        RECT 361.520 526.120 362.420 606.420 ;
        RECT 364.820 605.800 516.020 606.420 ;
        RECT 364.820 526.740 512.720 605.800 ;
        RECT 515.120 526.740 516.020 605.800 ;
        RECT 518.420 526.740 666.320 606.420 ;
        RECT 668.720 526.740 669.620 606.420 ;
        RECT 364.820 526.120 669.620 526.740 ;
        RECT 672.020 526.120 819.920 606.420 ;
        RECT 100.620 97.415 819.920 526.120 ;
        RECT 822.320 97.415 823.220 1105.505 ;
        RECT 825.620 1016.745 973.520 1105.505 ;
        RECT 975.920 1016.745 976.820 1105.505 ;
        RECT 979.220 1016.745 1127.120 1105.505 ;
        RECT 1129.520 1016.745 1130.420 1105.505 ;
        RECT 1132.820 1016.745 1280.720 1105.505 ;
        RECT 825.620 371.775 1280.720 1016.745 ;
        RECT 825.620 97.415 973.520 371.775 ;
        RECT 975.920 97.415 976.820 371.775 ;
        RECT 979.220 97.415 1127.120 371.775 ;
        RECT 1129.520 97.415 1130.420 371.775 ;
        RECT 1132.820 97.415 1280.720 371.775 ;
        RECT 1283.120 97.415 1284.020 1105.505 ;
        RECT 1286.420 97.415 1296.905 1105.505 ;
  END
END osiris_i_mem
END LIBRARY

